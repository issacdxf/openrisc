
//- 0-In CDC V2.5d (suse9_x86) 06/05/07

//-----------------------------------------------------------------
// CDC Control File
// Created Thu Sep 17 12:05:28 2009
//-----------------------------------------------------------------


module zin_cdc_ctrl_des_0;


`include "/export/home/user/wangyl/rtlqa_env/digital/impl/cdc/run_dir/0in_cdc_param.inc"


endmodule


