
module SNPS_CLOCK_GATE_OBS_tiny_des_round ( TE, net1780, hclk, test_se, 
        test_si, test_so );
  input TE, net1780, hclk, test_se, test_si;
  output test_so;
  wire   net1790, net1792;

  AN2 main_gate ( .I1(TE), .I2(hclk), .O(net1790) );
  ND2 nand_0_0 ( .I1(net1780), .I2(TE), .O(net1792) );
  QDFZS U1 ( .D(net1792), .TD(test_si), .SEL(test_se), .CK(net1790), .Q(
        test_so) );
endmodule


module POWERMODULE_HIGH_tiny_des_round_0 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1771;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2P main_gate ( .I1(net1771), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1771) );
endmodule


module tiny_des_round ( hclk, POR, hresetn, stall, encrypt_in, encrypt_shift, 
        decrypt_shift, key_in, din, dout, test_mode, test_se, test_si );
  input [4:0] encrypt_shift;
  input [4:0] decrypt_shift;
  input [63:0] key_in;
  input [63:0] din;
  output [63:0] dout;
  input hclk, POR, hresetn, stall, encrypt_in, test_mode, test_se, test_si;
  wire   N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754, N1755,
         N1756, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765,
         N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775,
         N1776, N1777, N1778, CLKGATING_hclk_POWERGATING_hclk_N1778_0_0,
         net1780, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1508, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1645, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n1, n2, n56, n57, n83, n84, n400,
         n401, n432, n433, n1373, n1440, n1507, n1509, n1585, n1644, n1646,
         n1738, n1739, n1740, n1800, n1801, n1802, n1817, n1960, n1961, n2005,
         n2006, n2181, n2280, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2557;

  OA22P U1142 ( .A1(n2506), .A2(n1659), .B1(n1660), .B2(n2500), .O(n247) );
  OA22P U1222 ( .A1(n2529), .A2(n1720), .B1(n1721), .B2(n2533), .O(n275) );
  OA2222 U1456 ( .A1(n1640), .A2(n1647), .B1(n1642), .B2(n1658), .C1(n2491), 
        .C2(n1890), .D1(n2486), .D2(n1891), .O(n1638) );
  OA2222 U1457 ( .A1(n1640), .A2(n1891), .B1(n1642), .B2(n1641), .C1(n2491), 
        .C2(n1643), .D1(n2486), .D2(n1645), .O(n1662) );
  OA2222 U1550 ( .A1(n1503), .A2(n1708), .B1(n1505), .B2(n1719), .C1(n2474), 
        .C2(n1952), .D1(n2469), .D2(n1953), .O(n1703) );
  OA2222 U1552 ( .A1(n1503), .A2(n1953), .B1(n1505), .B2(n1705), .C1(n2475), 
        .C2(n1706), .D1(n2469), .D2(n1707), .O(n1722) );
  OR3B2P U1659 ( .I1(n884), .B1(n321), .B2(n878), .O(n1312) );
  OA2222 U1725 ( .A1(n1503), .A2(n1777), .B1(n1505), .B2(n1776), .C1(n2474), 
        .C2(n1504), .D1(n2469), .D2(n1506), .O(n1781) );
  OA2222 U1793 ( .A1(n1503), .A2(n1778), .B1(n1505), .B2(n1777), .C1(n2475), 
        .C2(n1776), .D1(n2469), .D2(n1504), .O(n1501) );
  OA2222 U1794 ( .A1(n2098), .A2(n2462), .B1(n2099), .B2(n2458), .C1(n2100), 
        .C2(n2454), .D1(n2089), .D2(n2450), .O(n1504) );
  OA2222 U1795 ( .A1(n2102), .A2(n2462), .B1(n2103), .B2(n2458), .C1(n2104), 
        .C2(n2454), .D1(n2097), .D2(n2450), .O(n1776) );
  OA2222 U1796 ( .A1(n2107), .A2(n2462), .B1(n2108), .B2(n2458), .C1(n2109), 
        .C2(n2454), .D1(n2101), .D2(n2450), .O(n1777) );
  OA2222 U1798 ( .A1(n1503), .A2(n1506), .B1(n1505), .B2(n1508), .C1(n2475), 
        .C2(n1510), .D1(n2469), .D2(n1778), .O(n2053) );
  OA2222 U1799 ( .A1(n2111), .A2(n2462), .B1(n2112), .B2(n2458), .C1(n2113), 
        .C2(n2454), .D1(n2106), .D2(n2450), .O(n1778) );
  OA2222 U1800 ( .A1(n2115), .A2(n2462), .B1(n2116), .B2(n2458), .C1(n2117), 
        .C2(n2454), .D1(n2110), .D2(n2450), .O(n1510) );
  OA2222 U1801 ( .A1(n2119), .A2(n2462), .B1(n2120), .B2(n2458), .C1(n2121), 
        .C2(n2454), .D1(n2114), .D2(n2450), .O(n1508) );
  OA2222 U1802 ( .A1(n2091), .A2(n2462), .B1(n2093), .B2(n2458), .C1(n2095), 
        .C2(n2454), .D1(n2118), .D2(n2450), .O(n1506) );
  OA2222 U1996 ( .A1(n1640), .A2(n1890), .B1(n1642), .B2(n1891), .C1(n2491), 
        .C2(n1641), .D1(n2486), .D2(n1643), .O(n1657) );
  OA2222 U1997 ( .A1(n2446), .A2(n2223), .B1(n2442), .B2(n2224), .C1(n2438), 
        .C2(n2225), .D1(n2434), .D2(n2226), .O(n1643) );
  OA2222 U1998 ( .A1(n2446), .A2(n2227), .B1(n2442), .B2(n2228), .C1(n2438), 
        .C2(n2229), .D1(n2434), .D2(n2230), .O(n1641) );
  OA2222 U1999 ( .A1(n2446), .A2(n2231), .B1(n2442), .B2(n2232), .C1(n2438), 
        .C2(n2233), .D1(n2434), .D2(n2234), .O(n1891) );
  OA2222 U2002 ( .A1(n2446), .A2(n2236), .B1(n2442), .B2(n2237), .C1(n2438), 
        .C2(n2238), .D1(n2434), .D2(n2239), .O(n1645) );
  OA2222 U2003 ( .A1(n2446), .A2(n2240), .B1(n2442), .B2(n2241), .C1(n2438), 
        .C2(n2242), .D1(n2434), .D2(n2243), .O(n1647) );
  OA2222 U2005 ( .A1(n2446), .A2(n2244), .B1(n2442), .B2(n2245), .C1(n2438), 
        .C2(n2246), .D1(n2434), .D2(n2247), .O(n1658) );
  OA2222 U2007 ( .A1(n2446), .A2(n2248), .B1(n2442), .B2(n2249), .C1(n2438), 
        .C2(n2250), .D1(n2434), .D2(n2251), .O(n1890) );
  OA2222 U2107 ( .A1(n1503), .A2(n1952), .B1(n1505), .B2(n1953), .C1(n2474), 
        .C2(n1705), .D1(n2469), .D2(n1706), .O(n1718) );
  OA2222 U2108 ( .A1(n2462), .A2(n2223), .B1(n2458), .B2(n2224), .C1(n2454), 
        .C2(n2225), .D1(n2450), .D2(n2226), .O(n1706) );
  OA2222 U2109 ( .A1(n2462), .A2(n2227), .B1(n2458), .B2(n2228), .C1(n2454), 
        .C2(n2229), .D1(n2450), .D2(n2230), .O(n1705) );
  OA2222 U2110 ( .A1(n2462), .A2(n2231), .B1(n2458), .B2(n2232), .C1(n2454), 
        .C2(n2233), .D1(n2450), .D2(n2234), .O(n1953) );
  OA2222 U2113 ( .A1(n2462), .A2(n2236), .B1(n2458), .B2(n2237), .C1(n2454), 
        .C2(n2238), .D1(n2450), .D2(n2239), .O(n1707) );
  OA2222 U2114 ( .A1(n2462), .A2(n2240), .B1(n2458), .B2(n2241), .C1(n2454), 
        .C2(n2242), .D1(n2450), .D2(n2243), .O(n1708) );
  OA2222 U2116 ( .A1(n2462), .A2(n2244), .B1(n2458), .B2(n2245), .C1(n2454), 
        .C2(n2246), .D1(n2450), .D2(n2247), .O(n1719) );
  OA2222 U2118 ( .A1(n2462), .A2(n2248), .B1(n2458), .B2(n2249), .C1(n2454), 
        .C2(n2250), .D1(n2450), .D2(n2251), .O(n1952) );
  OAI222 U2179 ( .A1(n235), .A2(n236), .B1(n237), .B2(n238), .C1(n239), .C2(
        n240), .O(n234) );
  OAI222 U2180 ( .A1(n263), .A2(n2390), .B1(n265), .B2(n266), .C1(n267), .C2(
        n268), .O(n262) );
  OAI2222 U2181 ( .A1(n352), .A2(n353), .B1(n354), .B2(n355), .C1(n356), .C2(
        n357), .D1(n358), .D2(n359), .O(n346) );
  AOI2222 U2182 ( .A1(n911), .A2(n912), .B1(n513), .B2(n913), .C1(n914), .C2(
        n908), .D1(n915), .D2(n2325), .O(n905) );
  AOI2222 U2183 ( .A1(n931), .A2(n932), .B1(n2316), .B2(n933), .C1(n934), .C2(
        n928), .D1(n935), .D2(n468), .O(n925) );
  AOI2222 U2184 ( .A1(n2497), .A2(n1382), .B1(n2494), .B2(n1391), .C1(n2489), 
        .C2(n1392), .D1(n2484), .D2(n1393), .O(n1372) );
  AOI2222 U2185 ( .A1(n2481), .A2(n1449), .B1(n2477), .B2(n1457), .C1(n2472), 
        .C2(n1458), .D1(n2467), .D2(n1459), .O(n1439) );
  OAI2222 U2186 ( .A1(n1503), .A2(n1504), .B1(n1505), .B2(n1506), .C1(n2475), 
        .C2(n1508), .D1(n2470), .D2(n1510), .O(n1502) );
  AOI2222 U2187 ( .A1(n1588), .A2(n2483), .B1(n1589), .B2(n2489), .C1(n1590), 
        .C2(n2493), .D1(n1591), .D2(n2497), .O(n1586) );
  OAI2222 U2188 ( .A1(n1640), .A2(n1641), .B1(n1642), .B2(n1643), .C1(n2491), 
        .C2(n1645), .D1(n2486), .D2(n1647), .O(n1639) );
  AOI2222 U2189 ( .A1(n2497), .A2(n1651), .B1(n2493), .B2(n1652), .C1(n2488), 
        .C2(n1653), .D1(n2483), .D2(n1654), .O(n1400) );
  AOI2222 U2190 ( .A1(n2481), .A2(n1697), .B1(n2476), .B2(n1698), .C1(n2471), 
        .C2(n1699), .D1(n2466), .D2(n1700), .O(n1469) );
  OAI2222 U2191 ( .A1(n1503), .A2(n1705), .B1(n1505), .B2(n1706), .C1(n2475), 
        .C2(n1707), .D1(n2470), .D2(n1708), .O(n1704) );
  AOI2222 U2192 ( .A1(n2481), .A2(n1712), .B1(n2476), .B2(n1713), .C1(n2471), 
        .C2(n1714), .D1(n2466), .D2(n1715), .O(n1464) );
  NR6 U2193 ( .I1(n1730), .I2(n1731), .I3(n949), .I4(n79), .I5(n55), .I6(n947), 
        .O(n1729) );
  AOI2222 U2194 ( .A1(n2481), .A2(n1758), .B1(n2476), .B2(n1759), .C1(n2471), 
        .C2(n1760), .D1(n2466), .D2(n1761), .O(n1523) );
  AOI2222 U2195 ( .A1(n1765), .A2(n2466), .B1(n1535), .B2(n2473), .C1(n1534), 
        .C2(n2476), .D1(n1533), .D2(n2481), .O(n1763) );
  AOI2222 U2196 ( .A1(n2481), .A2(n1761), .B1(n2476), .B2(n1770), .C1(n2471), 
        .C2(n1771), .D1(n2466), .D2(n1772), .O(n1757) );
  OAI2222 U2197 ( .A1(n1503), .A2(n1508), .B1(n1505), .B2(n1510), .C1(n2475), 
        .C2(n1778), .D1(n2470), .D2(n1777), .O(n1782) );
  AOI2222 U2198 ( .A1(n2481), .A2(n1785), .B1(n2476), .B2(n1786), .C1(n2471), 
        .C2(n1787), .D1(n2466), .D2(n1788), .O(n1520) );
  NR6 U2199 ( .I1(n1792), .I2(n1793), .I3(n981), .I4(n106), .I5(n82), .I6(n979), .O(n1791) );
  AOI2222 U2200 ( .A1(n2497), .A2(n1819), .B1(n2493), .B2(n1820), .C1(n2488), 
        .C2(n1821), .D1(n2483), .D2(n1822), .O(n1581) );
  AOI2222 U2201 ( .A1(n1826), .A2(n2483), .B1(n1588), .B2(n2489), .C1(n1589), 
        .C2(n2493), .D1(n1590), .D2(n2497), .O(n1824) );
  AOI2222 U2202 ( .A1(n2497), .A2(n1822), .B1(n2493), .B2(n1829), .C1(n2488), 
        .C2(n1830), .D1(n2483), .D2(n1831), .O(n1818) );
  AOI2222 U2203 ( .A1(n1574), .A2(n2483), .B1(n1573), .B2(n2489), .C1(n1572), 
        .C2(n2493), .D1(n1835), .D2(n2497), .O(n1834) );
  AOI2222 U2204 ( .A1(n1835), .A2(n2483), .B1(n1836), .B2(n2489), .C1(n1837), 
        .C2(n2493), .D1(n1575), .D2(n2497), .O(n1833) );
  AOI2222 U2205 ( .A1(n2497), .A2(n1635), .B1(n2493), .B2(n1886), .C1(n2488), 
        .C2(n1887), .D1(n2483), .D2(n1888), .O(n1404) );
  AOI2222 U2206 ( .A1(n2497), .A2(n1894), .B1(n2493), .B2(n1651), .C1(n2488), 
        .C2(n1652), .D1(n2483), .D2(n1653), .O(n1883) );
  AOI2222 U2207 ( .A1(n2497), .A2(n1886), .B1(n2493), .B2(n1887), .C1(n2488), 
        .C2(n1888), .D1(n2483), .D2(n1632), .O(n1631) );
  AOI2222 U2208 ( .A1(n2481), .A2(n1700), .B1(n2476), .B2(n1940), .C1(n2471), 
        .C2(n1941), .D1(n2466), .D2(n1942), .O(n1468) );
  AOI2222 U2209 ( .A1(n2481), .A2(n1940), .B1(n2476), .B2(n1941), .C1(n2471), 
        .C2(n1942), .D1(n2466), .D2(n1697), .O(n1701) );
  AOI2222 U2210 ( .A1(n2480), .A2(n1698), .B1(n2476), .B2(n1699), .C1(n2471), 
        .C2(n1700), .D1(n2466), .D2(n1940), .O(n1725) );
  AOI2222 U2211 ( .A1(n2480), .A2(n1947), .B1(n2476), .B2(n1712), .C1(n2471), 
        .C2(n1713), .D1(n2466), .D2(n1714), .O(n1936) );
  AOI2222 U2212 ( .A1(n2480), .A2(n1715), .B1(n2477), .B2(n1948), .C1(n2471), 
        .C2(n1949), .D1(n2467), .D2(n1947), .O(n1711) );
  AOI2222 U2213 ( .A1(n2497), .A2(n1845), .B1(n2494), .B2(n1846), .C1(n2488), 
        .C2(n1990), .D1(n2484), .D2(n1991), .O(n1584) );
  AOI2222 U2214 ( .A1(n2497), .A2(n1821), .B1(n2494), .B2(n1822), .C1(n2488), 
        .C2(n1829), .D1(n2484), .D2(n1830), .O(n1567) );
  AOI2222 U2215 ( .A1(n2497), .A2(n1846), .B1(n2494), .B2(n1990), .C1(n2488), 
        .C2(n1991), .D1(n2484), .D2(n1995), .O(n1577) );
  AOI2222 U2216 ( .A1(n2497), .A2(n1836), .B1(n2494), .B2(n1835), .C1(n2488), 
        .C2(n1572), .D1(n2484), .D2(n1573), .O(n1839) );
  AOI2222 U2217 ( .A1(n2480), .A2(n1771), .B1(n2477), .B2(n1772), .C1(n2472), 
        .C2(n1758), .D1(n2467), .D2(n1759), .O(n1513) );
  AOI2222 U2218 ( .A1(n2480), .A2(n1787), .B1(n2477), .B2(n1788), .C1(n2472), 
        .C2(n2041), .D1(n2467), .D2(n2042), .O(n1527) );
  AOI2222 U2219 ( .A1(n2480), .A2(n2045), .B1(n2477), .B2(n1785), .C1(n2472), 
        .C2(n1786), .D1(n2467), .D2(n1787), .O(n1528) );
  AOI2222 U2220 ( .A1(n2480), .A2(n1788), .B1(n2477), .B2(n2041), .C1(n2472), 
        .C2(n2042), .D1(n2467), .D2(n2045), .O(n1518) );
  AOI2222 U2221 ( .A1(n2480), .A2(n1760), .B1(n2477), .B2(n1761), .C1(n2472), 
        .C2(n1770), .D1(n2467), .D2(n1771), .O(n1515) );
  AOI2222 U2222 ( .A1(n2480), .A2(n1772), .B1(n2477), .B2(n1758), .C1(n2472), 
        .C2(n1759), .D1(n2467), .D2(n1760), .O(n1768) );
  AOI2222 U2223 ( .A1(n2480), .A2(n2041), .B1(n2477), .B2(n2042), .C1(n2472), 
        .C2(n2045), .D1(n2467), .D2(n1785), .O(n1790) );
  AOI2222 U2224 ( .A1(n2480), .A2(n1770), .B1(n2477), .B2(n1771), .C1(n2472), 
        .C2(n1772), .D1(n2467), .D2(n1758), .O(n1524) );
  OAI2222 U2225 ( .A1(n2089), .A2(n2465), .B1(n2091), .B2(n2460), .C1(n2093), 
        .C2(n2457), .D1(n2095), .D2(n2452), .O(n1758) );
  OAI2222 U2226 ( .A1(n2097), .A2(n2465), .B1(n2098), .B2(n2458), .C1(n2099), 
        .C2(n2457), .D1(n2100), .D2(n2450), .O(n1772) );
  OAI2222 U2227 ( .A1(n2101), .A2(n2465), .B1(n2102), .B2(n2458), .C1(n2103), 
        .C2(n2457), .D1(n2104), .D2(n2450), .O(n1771) );
  AOI2222 U2228 ( .A1(n2480), .A2(n1759), .B1(n2477), .B2(n1760), .C1(n2472), 
        .C2(n1761), .D1(n2467), .D2(n1770), .O(n2036) );
  OAI2222 U2229 ( .A1(n2106), .A2(n2465), .B1(n2107), .B2(n2459), .C1(n2108), 
        .C2(n2457), .D1(n2109), .D2(n2451), .O(n1770) );
  OAI2222 U2230 ( .A1(n2110), .A2(n2465), .B1(n2111), .B2(n2459), .C1(n2112), 
        .C2(n2457), .D1(n2113), .D2(n2451), .O(n1761) );
  OAI2222 U2231 ( .A1(n2114), .A2(n2465), .B1(n2115), .B2(n2459), .C1(n2116), 
        .C2(n2457), .D1(n2117), .D2(n2451), .O(n1760) );
  OAI2222 U2232 ( .A1(n2118), .A2(n2465), .B1(n2119), .B2(n2459), .C1(n2120), 
        .C2(n2457), .D1(n2121), .D2(n2451), .O(n1759) );
  AOI2222 U2233 ( .A1(n2480), .A2(n1786), .B1(n2477), .B2(n1787), .C1(n2472), 
        .C2(n1788), .D1(n2467), .D2(n2041), .O(n2050) );
  OAI2222 U2234 ( .A1(n2113), .A2(n2465), .B1(n2106), .B2(n2459), .C1(n2107), 
        .C2(n2457), .D1(n2108), .D2(n2451), .O(n2041) );
  OAI2222 U2235 ( .A1(n2117), .A2(n2464), .B1(n2110), .B2(n2459), .C1(n2111), 
        .C2(n2456), .D1(n2112), .D2(n2451), .O(n1788) );
  OAI2222 U2236 ( .A1(n2121), .A2(n2464), .B1(n2114), .B2(n2459), .C1(n2115), 
        .C2(n2456), .D1(n2116), .D2(n2451), .O(n1787) );
  AOI2222 U2237 ( .A1(n2480), .A2(n2042), .B1(n2477), .B2(n2045), .C1(n2472), 
        .C2(n1785), .D1(n2467), .D2(n1786), .O(n2040) );
  OAI2222 U2238 ( .A1(n2095), .A2(n2464), .B1(n2118), .B2(n2459), .C1(n2119), 
        .C2(n2456), .D1(n2120), .D2(n2451), .O(n1786) );
  OAI2222 U2239 ( .A1(n2100), .A2(n2464), .B1(n2089), .B2(n2459), .C1(n2091), 
        .C2(n2456), .D1(n2093), .D2(n2451), .O(n1785) );
  OAI2222 U2240 ( .A1(n2104), .A2(n2464), .B1(n2097), .B2(n2459), .C1(n2098), 
        .C2(n2456), .D1(n2099), .D2(n2451), .O(n2045) );
  OAI2222 U2241 ( .A1(n2109), .A2(n2464), .B1(n2101), .B2(n2459), .C1(n2102), 
        .C2(n2456), .D1(n2103), .D2(n2451), .O(n2042) );
  AOI2222 U2242 ( .A1(n2480), .A2(n2133), .B1(n2477), .B2(n1532), .C1(n2472), 
        .C2(n1533), .D1(n2467), .D2(n1534), .O(n2129) );
  AOI2222 U2243 ( .A1(n2480), .A2(n1535), .B1(n2477), .B2(n1765), .C1(n2472), 
        .C2(n2134), .D1(n2467), .D2(n2133), .O(n1530) );
  AOI2222 U2244 ( .A1(n2479), .A2(n1534), .B1(n2477), .B2(n1535), .C1(n2472), 
        .C2(n1765), .D1(n2467), .D2(n2134), .O(n2130) );
  OAI2222 U2245 ( .A1(n2108), .A2(n2464), .B1(n2109), .B2(n2459), .C1(n2101), 
        .C2(n2456), .D1(n2102), .D2(n2451), .O(n1765) );
  OAI2222 U2246 ( .A1(n2112), .A2(n2464), .B1(n2113), .B2(n2459), .C1(n2106), 
        .C2(n2456), .D1(n2107), .D2(n2451), .O(n1535) );
  OAI2222 U2247 ( .A1(n2116), .A2(n2464), .B1(n2117), .B2(n2459), .C1(n2110), 
        .C2(n2456), .D1(n2111), .D2(n2451), .O(n1534) );
  AOI2222 U2248 ( .A1(n2479), .A2(n2134), .B1(n2478), .B2(n2133), .C1(n2472), 
        .C2(n1532), .D1(n2468), .D2(n1533), .O(n1764) );
  OAI2222 U2249 ( .A1(n2120), .A2(n2464), .B1(n2121), .B2(n2459), .C1(n2114), 
        .C2(n2456), .D1(n2115), .D2(n2451), .O(n1533) );
  OAI2222 U2250 ( .A1(n2093), .A2(n2464), .B1(n2095), .B2(n2459), .C1(n2118), 
        .C2(n2456), .D1(n2119), .D2(n2451), .O(n1532) );
  OAI2222 U2251 ( .A1(n2099), .A2(n2464), .B1(n2100), .B2(n2460), .C1(n2089), 
        .C2(n2456), .D1(n2091), .D2(n2452), .O(n2133) );
  OAI2222 U2252 ( .A1(n2103), .A2(n2464), .B1(n2104), .B2(n2460), .C1(n2097), 
        .C2(n2456), .D1(n2098), .D2(n2452), .O(n2134) );
  AOI2222 U2253 ( .A1(n2497), .A2(n1820), .B1(n2494), .B2(n1821), .C1(n2489), 
        .C2(n1822), .D1(n2484), .D2(n1829), .O(n2003) );
  OAI2222 U2254 ( .A1(n2110), .A2(n2449), .B1(n2111), .B2(n2442), .C1(n2112), 
        .C2(n2441), .D1(n2437), .D2(n2113), .O(n1822) );
  OAI2222 U2255 ( .A1(n2446), .A2(n2114), .B1(n2442), .B2(n2115), .C1(n2441), 
        .C2(n2116), .D1(n2437), .D2(n2117), .O(n1821) );
  OAI2222 U2256 ( .A1(n2446), .A2(n2118), .B1(n2442), .B2(n2119), .C1(n2441), 
        .C2(n2120), .D1(n2437), .D2(n2121), .O(n1820) );
  OAI2222 U2257 ( .A1(n2446), .A2(n2089), .B1(n2442), .B2(n2091), .C1(n2441), 
        .C2(n2093), .D1(n2437), .D2(n2095), .O(n1819) );
  OAI2222 U2258 ( .A1(n2446), .A2(n2097), .B1(n2442), .B2(n2098), .C1(n2441), 
        .C2(n2099), .D1(n2437), .D2(n2100), .O(n1831) );
  OAI2222 U2259 ( .A1(n2446), .A2(n2101), .B1(n2442), .B2(n2102), .C1(n2441), 
        .C2(n2103), .D1(n2437), .D2(n2104), .O(n1830) );
  OAI2222 U2260 ( .A1(n2446), .A2(n2106), .B1(n2442), .B2(n2107), .C1(n2441), 
        .C2(n2108), .D1(n2437), .D2(n2109), .O(n1829) );
  AOI2222 U2261 ( .A1(n2496), .A2(n1844), .B1(n2494), .B2(n1845), .C1(n2489), 
        .C2(n1846), .D1(n2484), .D2(n1990), .O(n1998) );
  OAI2222 U2262 ( .A1(n2446), .A2(n2113), .B1(n2443), .B2(n2106), .C1(n2441), 
        .C2(n2107), .D1(n2437), .D2(n2108), .O(n1990) );
  OAI2222 U2263 ( .A1(n2446), .A2(n2117), .B1(n2443), .B2(n2110), .C1(n2440), 
        .C2(n2111), .D1(n2436), .D2(n2112), .O(n1846) );
  OAI2222 U2264 ( .A1(n2447), .A2(n2121), .B1(n2443), .B2(n2114), .C1(n2440), 
        .C2(n2115), .D1(n2436), .D2(n2116), .O(n1845) );
  OAI2222 U2265 ( .A1(n2447), .A2(n2095), .B1(n2443), .B2(n2118), .C1(n2440), 
        .C2(n2119), .D1(n2436), .D2(n2120), .O(n1844) );
  OAI2222 U2266 ( .A1(n2447), .A2(n2100), .B1(n2443), .B2(n2089), .C1(n2440), 
        .C2(n2091), .D1(n2436), .D2(n2093), .O(n1843) );
  OAI2222 U2267 ( .A1(n2447), .A2(n2104), .B1(n2443), .B2(n2097), .C1(n2440), 
        .C2(n2098), .D1(n2436), .D2(n2099), .O(n1995) );
  OAI2222 U2268 ( .A1(n2447), .A2(n2109), .B1(n2443), .B2(n2101), .C1(n2440), 
        .C2(n2102), .D1(n2436), .D2(n2103), .O(n1991) );
  AOI2222 U2269 ( .A1(n2496), .A2(n1837), .B1(n2494), .B2(n1836), .C1(n2489), 
        .C2(n1835), .D1(n2484), .D2(n1572), .O(n1570) );
  OAI2222 U2270 ( .A1(n2447), .A2(n2098), .B1(n2443), .B2(n2099), .C1(n2440), 
        .C2(n2100), .D1(n2436), .D2(n2089), .O(n1572) );
  OAI2222 U2271 ( .A1(n2447), .A2(n2102), .B1(n2443), .B2(n2103), .C1(n2440), 
        .C2(n2104), .D1(n2436), .D2(n2097), .O(n1835) );
  OAI2222 U2272 ( .A1(n2447), .A2(n2107), .B1(n2443), .B2(n2108), .C1(n2440), 
        .C2(n2109), .D1(n2436), .D2(n2101), .O(n1836) );
  OAI2222 U2273 ( .A1(n2111), .A2(n2449), .B1(n2112), .B2(n2442), .C1(n2440), 
        .C2(n2113), .D1(n2436), .D2(n2106), .O(n1837) );
  OAI2222 U2274 ( .A1(n2447), .A2(n2115), .B1(n2443), .B2(n2116), .C1(n2440), 
        .C2(n2117), .D1(n2436), .D2(n2110), .O(n1575) );
  OAI2222 U2275 ( .A1(n2447), .A2(n2119), .B1(n2443), .B2(n2120), .C1(n2440), 
        .C2(n2121), .D1(n2436), .D2(n2114), .O(n1574) );
  OAI2222 U2276 ( .A1(n2447), .A2(n2091), .B1(n2443), .B2(n2093), .C1(n2440), 
        .C2(n2095), .D1(n2436), .D2(n2118), .O(n1573) );
  AOI2222 U2277 ( .A1(n2496), .A2(n1588), .B1(n2494), .B2(n1826), .C1(n2489), 
        .C2(n2179), .D1(n2484), .D2(n2180), .O(n1587) );
  AOI2222 U2278 ( .A1(n2496), .A2(n2179), .B1(n2494), .B2(n2180), .C1(n2489), 
        .C2(n1591), .D1(n2484), .D2(n1590), .O(n1825) );
  OAI2222 U2279 ( .A1(n2447), .A2(n2120), .B1(n2443), .B2(n2121), .C1(n2440), 
        .C2(n2114), .D1(n2436), .D2(n2115), .O(n1590) );
  OAI2222 U2280 ( .A1(n2447), .A2(n2093), .B1(n2443), .B2(n2095), .C1(n2440), 
        .C2(n2118), .D1(n2436), .D2(n2119), .O(n1591) );
  OAI2222 U2281 ( .A1(n2447), .A2(n2099), .B1(n2443), .B2(n2100), .C1(n2440), 
        .C2(n2089), .D1(n2436), .D2(n2091), .O(n2180) );
  AOI2222 U2282 ( .A1(n2496), .A2(n1589), .B1(n2494), .B2(n1588), .C1(n2489), 
        .C2(n1826), .D1(n2484), .D2(n2179), .O(n2177) );
  OAI2222 U2283 ( .A1(n2447), .A2(n2103), .B1(n2444), .B2(n2104), .C1(n2439), 
        .C2(n2097), .D1(n2435), .D2(n2098), .O(n2179) );
  OAI2222 U2284 ( .A1(n2447), .A2(n2108), .B1(n2444), .B2(n2109), .C1(n2439), 
        .C2(n2101), .D1(n2435), .D2(n2102), .O(n1826) );
  OAI2222 U2285 ( .A1(n2112), .A2(n2449), .B1(n2444), .B2(n2113), .C1(n2439), 
        .C2(n2106), .D1(n2435), .D2(n2107), .O(n1588) );
  OAI2222 U2286 ( .A1(n2448), .A2(n2116), .B1(n2444), .B2(n2117), .C1(n2439), 
        .C2(n2110), .D1(n2435), .D2(n2111), .O(n1589) );
  OAI222 U2287 ( .A1(n2190), .A2(n637), .B1(n2196), .B2(n2198), .C1(n2199), 
        .C2(n2193), .O(n2197) );
  AOI2222 U2288 ( .A1(n2496), .A2(n1887), .B1(n2494), .B2(n1888), .C1(n2489), 
        .C2(n1632), .D1(n2484), .D2(n1633), .O(n1626) );
  AOI2222 U2289 ( .A1(n2496), .A2(n1392), .B1(n2494), .B2(n1393), .C1(n2489), 
        .C2(n1376), .D1(n2484), .D2(n1378), .O(n1900) );
  OAI2222 U2290 ( .A1(n2448), .A2(n2239), .B1(n2444), .B2(n2240), .C1(n2439), 
        .C2(n2241), .D1(n2435), .D2(n2242), .O(n1376) );
  OAI2222 U2291 ( .A1(n2448), .A2(n2226), .B1(n2444), .B2(n2236), .C1(n2439), 
        .C2(n2237), .D1(n2435), .D2(n2238), .O(n1393) );
  OAI2222 U2292 ( .A1(n2448), .A2(n2230), .B1(n2444), .B2(n2223), .C1(n2439), 
        .C2(n2224), .D1(n2435), .D2(n2225), .O(n1392) );
  AOI2222 U2293 ( .A1(n2496), .A2(n1378), .B1(n2494), .B2(n1380), .C1(n2489), 
        .C2(n1382), .D1(n2484), .D2(n1391), .O(n1389) );
  OAI2222 U2294 ( .A1(n2448), .A2(n2234), .B1(n2444), .B2(n2227), .C1(n2439), 
        .C2(n2228), .D1(n2435), .D2(n2229), .O(n1391) );
  OAI2222 U2295 ( .A1(n2448), .A2(n2251), .B1(n2444), .B2(n2231), .C1(n2439), 
        .C2(n2232), .D1(n2435), .D2(n2233), .O(n1382) );
  OAI2222 U2296 ( .A1(n2448), .A2(n2247), .B1(n2444), .B2(n2248), .C1(n2439), 
        .C2(n2249), .D1(n2435), .D2(n2250), .O(n1380) );
  OAI2222 U2297 ( .A1(n2448), .A2(n2243), .B1(n2444), .B2(n2244), .C1(n2439), 
        .C2(n2245), .D1(n2435), .D2(n2246), .O(n1378) );
  AOI2222 U2298 ( .A1(n2496), .A2(n1634), .B1(n2494), .B2(n1635), .C1(n2489), 
        .C2(n1886), .D1(n2484), .D2(n1887), .O(n2221) );
  OAI2222 U2299 ( .A1(n2448), .A2(n2238), .B1(n2444), .B2(n2239), .C1(n2439), 
        .C2(n2240), .D1(n2435), .D2(n2241), .O(n1887) );
  OAI2222 U2300 ( .A1(n2448), .A2(n2225), .B1(n2444), .B2(n2226), .C1(n2439), 
        .C2(n2236), .D1(n2435), .D2(n2237), .O(n1886) );
  OAI2222 U2301 ( .A1(n2448), .A2(n2229), .B1(n2444), .B2(n2230), .C1(n2439), 
        .C2(n2223), .D1(n2435), .D2(n2224), .O(n1635) );
  OAI2222 U2302 ( .A1(n2448), .A2(n2233), .B1(n2444), .B2(n2234), .C1(n2439), 
        .C2(n2227), .D1(n2435), .D2(n2228), .O(n1634) );
  OAI2222 U2303 ( .A1(n2448), .A2(n2250), .B1(n2444), .B2(n2251), .C1(n2439), 
        .C2(n2231), .D1(n2435), .D2(n2232), .O(n1633) );
  OAI2222 U2304 ( .A1(n2448), .A2(n2246), .B1(n2445), .B2(n2247), .C1(n2438), 
        .C2(n2248), .D1(n2434), .D2(n2249), .O(n1632) );
  OAI2222 U2305 ( .A1(n2448), .A2(n2242), .B1(n2445), .B2(n2243), .C1(n2438), 
        .C2(n2244), .D1(n2434), .D2(n2245), .O(n1888) );
  AOI2222 U2306 ( .A1(n2496), .A2(n1896), .B1(n2494), .B2(n1894), .C1(n2489), 
        .C2(n1651), .D1(n2484), .D2(n1652), .O(n1386) );
  AOI2222 U2307 ( .A1(n2496), .A2(n1895), .B1(n2493), .B2(n1896), .C1(n2488), 
        .C2(n1894), .D1(n2483), .D2(n1651), .O(n1399) );
  OAI2222 U2308 ( .A1(n2449), .A2(n2241), .B1(n2445), .B2(n2242), .C1(n2438), 
        .C2(n2243), .D1(n2434), .D2(n2244), .O(n1651) );
  OAI2222 U2309 ( .A1(n2448), .A2(n2237), .B1(n2445), .B2(n2238), .C1(n2438), 
        .C2(n2239), .D1(n2434), .D2(n2240), .O(n1894) );
  OAI2222 U2310 ( .A1(n2449), .A2(n2224), .B1(n2445), .B2(n2225), .C1(n2438), 
        .C2(n2226), .D1(n2434), .D2(n2236), .O(n1896) );
  OAI2222 U2311 ( .A1(n2449), .A2(n2228), .B1(n2445), .B2(n2229), .C1(n2438), 
        .C2(n2230), .D1(n2434), .D2(n2223), .O(n1895) );
  OAI2222 U2312 ( .A1(n2449), .A2(n2232), .B1(n2445), .B2(n2233), .C1(n2438), 
        .C2(n2234), .D1(n2434), .D2(n2227), .O(n1654) );
  OAI2222 U2313 ( .A1(n2449), .A2(n2249), .B1(n2445), .B2(n2250), .C1(n2438), 
        .C2(n2251), .D1(n2434), .D2(n2231), .O(n1653) );
  OAI2222 U2314 ( .A1(n2446), .A2(n2245), .B1(n2442), .B2(n2246), .C1(n2438), 
        .C2(n2247), .D1(n2434), .D2(n2248), .O(n1652) );
  OAI222 U2315 ( .A1(n2267), .A2(n658), .B1(n2273), .B2(n2274), .C1(n2275), 
        .C2(n2270), .O(n2272) );
  AOI2222 U2316 ( .A1(n2479), .A2(n1941), .B1(n2478), .B2(n1942), .C1(n2473), 
        .C2(n1697), .D1(n2468), .D2(n1698), .O(n1726) );
  AOI2222 U2317 ( .A1(n2479), .A2(n1445), .B1(n2478), .B2(n1447), .C1(n2473), 
        .C2(n1449), .D1(n2468), .D2(n1457), .O(n1455) );
  OAI2222 U2318 ( .A1(n2464), .A2(n2234), .B1(n2460), .B2(n2227), .C1(n2456), 
        .C2(n2228), .D1(n2452), .D2(n2229), .O(n1457) );
  OAI2222 U2319 ( .A1(n2464), .A2(n2251), .B1(n2460), .B2(n2231), .C1(n2456), 
        .C2(n2232), .D1(n2452), .D2(n2233), .O(n1449) );
  OAI2222 U2320 ( .A1(n2464), .A2(n2247), .B1(n2460), .B2(n2248), .C1(n2456), 
        .C2(n2249), .D1(n2452), .D2(n2250), .O(n1447) );
  AOI2222 U2321 ( .A1(n2479), .A2(n1458), .B1(n2478), .B2(n1459), .C1(n2473), 
        .C2(n1443), .D1(n2468), .D2(n1445), .O(n1955) );
  OAI2222 U2322 ( .A1(n2463), .A2(n2243), .B1(n2460), .B2(n2244), .C1(n2455), 
        .C2(n2245), .D1(n2452), .D2(n2246), .O(n1445) );
  OAI2222 U2323 ( .A1(n2463), .A2(n2239), .B1(n2460), .B2(n2240), .C1(n2455), 
        .C2(n2241), .D1(n2452), .D2(n2242), .O(n1443) );
  OAI2222 U2324 ( .A1(n2463), .A2(n2226), .B1(n2460), .B2(n2236), .C1(n2455), 
        .C2(n2237), .D1(n2452), .D2(n2238), .O(n1459) );
  OAI2222 U2325 ( .A1(n2463), .A2(n2230), .B1(n2460), .B2(n2223), .C1(n2455), 
        .C2(n2224), .D1(n2452), .D2(n2225), .O(n1458) );
  AOI2222 U2326 ( .A1(n2479), .A2(n1699), .B1(n2478), .B2(n1700), .C1(n2473), 
        .C2(n1940), .D1(n2468), .D2(n1941), .O(n2299) );
  OAI2222 U2327 ( .A1(n2463), .A2(n2238), .B1(n2460), .B2(n2239), .C1(n2455), 
        .C2(n2240), .D1(n2452), .D2(n2241), .O(n1941) );
  OAI2222 U2328 ( .A1(n2463), .A2(n2225), .B1(n2460), .B2(n2226), .C1(n2455), 
        .C2(n2236), .D1(n2452), .D2(n2237), .O(n1940) );
  OAI2222 U2329 ( .A1(n2463), .A2(n2229), .B1(n2460), .B2(n2230), .C1(n2455), 
        .C2(n2223), .D1(n2452), .D2(n2224), .O(n1700) );
  AOI2222 U2330 ( .A1(n2479), .A2(n1942), .B1(n2478), .B2(n1697), .C1(n2473), 
        .C2(n1698), .D1(n2468), .D2(n1699), .O(n1939) );
  OAI2222 U2331 ( .A1(n2463), .A2(n2233), .B1(n2460), .B2(n2234), .C1(n2455), 
        .C2(n2227), .D1(n2452), .D2(n2228), .O(n1699) );
  OAI2222 U2332 ( .A1(n2463), .A2(n2250), .B1(n2460), .B2(n2251), .C1(n2455), 
        .C2(n2231), .D1(n2452), .D2(n2232), .O(n1698) );
  OAI2222 U2333 ( .A1(n2463), .A2(n2246), .B1(n2460), .B2(n2247), .C1(n2455), 
        .C2(n2248), .D1(n2452), .D2(n2249), .O(n1697) );
  OAI2222 U2334 ( .A1(n2463), .A2(n2242), .B1(n2461), .B2(n2243), .C1(n2455), 
        .C2(n2244), .D1(n2453), .D2(n2245), .O(n1942) );
  AOI2222 U2335 ( .A1(n2479), .A2(n1949), .B1(n2478), .B2(n1947), .C1(n2473), 
        .C2(n1712), .D1(n2468), .D2(n1713), .O(n1453) );
  AOI2222 U2336 ( .A1(n2479), .A2(n1714), .B1(n2478), .B2(n1715), .C1(n2473), 
        .C2(n1948), .D1(n2468), .D2(n1949), .O(n1935) );
  AOI2222 U2337 ( .A1(n2479), .A2(n1948), .B1(n2478), .B2(n1949), .C1(n2473), 
        .C2(n1947), .D1(n2468), .D2(n1712), .O(n1465) );
  OAI2222 U2338 ( .A1(n2463), .A2(n2241), .B1(n2461), .B2(n2242), .C1(n2455), 
        .C2(n2243), .D1(n2453), .D2(n2244), .O(n1712) );
  OAI2222 U2339 ( .A1(n2463), .A2(n2237), .B1(n2461), .B2(n2238), .C1(n2455), 
        .C2(n2239), .D1(n2453), .D2(n2240), .O(n1947) );
  OAI2222 U2340 ( .A1(n2463), .A2(n2224), .B1(n2461), .B2(n2225), .C1(n2455), 
        .C2(n2226), .D1(n2453), .D2(n2236), .O(n1949) );
  AOI2222 U2341 ( .A1(n2479), .A2(n1713), .B1(n2476), .B2(n1714), .C1(n2471), 
        .C2(n1715), .D1(n2466), .D2(n1948), .O(n1452) );
  OAI2222 U2342 ( .A1(n2463), .A2(n2228), .B1(n2461), .B2(n2229), .C1(n2455), 
        .C2(n2230), .D1(n2453), .D2(n2223), .O(n1948) );
  OAI2222 U2343 ( .A1(n2463), .A2(n2232), .B1(n2461), .B2(n2233), .C1(n2455), 
        .C2(n2234), .D1(n2453), .D2(n2227), .O(n1715) );
  OAI2222 U2344 ( .A1(n2462), .A2(n2249), .B1(n2461), .B2(n2250), .C1(n2454), 
        .C2(n2251), .D1(n2453), .D2(n2231), .O(n1714) );
  OAI2222 U2345 ( .A1(n2462), .A2(n2245), .B1(n2461), .B2(n2246), .C1(n2454), 
        .C2(n2247), .D1(n2453), .D2(n2248), .O(n1713) );
  POWERMODULE_HIGH_tiny_des_round_0 POWERGATING_hclk_N1778_0 ( .CLK(hclk), 
        .EN(N1778), .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .TE(
        n2555), .ENOBS(net1780) );
  SNPS_CLOCK_GATE_OBS_tiny_des_round clk_gate_obs ( .TE(n2555), .net1780(
        net1780), .hclk(hclk), .test_se(test_se), .test_si(test_si), .test_so(
        n2557) );
  ND2 U2 ( .I1(n525), .I2(n1547), .O(n541) );
  BUF1 U3 ( .I(n458), .O(n2403) );
  NR2P U4 ( .I1(n613), .I2(n1912), .O(n224) );
  NR2T U5 ( .I1(n484), .I2(n483), .O(n932) );
  NR2T U6 ( .I1(n916), .I2(n511), .O(n912) );
  NR2T U7 ( .I1(n354), .I2(n634), .O(n2200) );
  NR2P U8 ( .I1(n1740), .I2(n374), .O(n650) );
  NR2T U9 ( .I1(n378), .I2(n655), .O(n2276) );
  INV2 U10 ( .I(n337), .O(n897) );
  XOR2P U11 ( .I1(n1636), .I2(n1637), .O(n254) );
  NR2T U12 ( .I1(n837), .I2(n275), .O(n842) );
  XOR2P U13 ( .I1(n1702), .I2(n1637), .O(n282) );
  XOR2 U14 ( .I1(n1884), .I2(n1388), .O(n186) );
  NR2P U15 ( .I1(n424), .I2(n2422), .O(n129) );
  NR2T U16 ( .I1(n2403), .I2(n774), .O(n1423) );
  INV3 U17 ( .I(n1002), .O(n101) );
  XOR2P U18 ( .I1(n1500), .I2(n1402), .O(n21) );
  XOR2P U19 ( .I1(n1569), .I2(n1402), .O(n44) );
  ND3P U20 ( .I1(n539), .I2(n40), .I3(n2396), .O(n37) );
  INV2 U21 ( .I(n868), .O(n1963) );
  XNR2P U22 ( .I1(n1371), .I2(din[14]), .O(n424) );
  NR2T U23 ( .I1(n22), .I2(n548), .O(n1107) );
  NR2P U24 ( .I1(n45), .I2(n525), .O(n1078) );
  INV3 U25 ( .I(n1041), .O(n215) );
  XOR2P U26 ( .I1(n2168), .I2(n2105), .O(n485) );
  XOR2P U27 ( .I1(n2001), .I2(n2002), .O(n850) );
  XOR2P U28 ( .I1(n1999), .I2(n1519), .O(n867) );
  XOR2P U29 ( .I1(n1993), .I2(n1994), .O(n309) );
  BUF1 U30 ( .I(n889), .O(n2335) );
  ND3 U31 ( .I1(n341), .I2(n319), .I3(n1321), .O(n895) );
  XOR2P U32 ( .I1(n1629), .I2(n1630), .O(n252) );
  INV3 U33 ( .I(n186), .O(n582) );
  INV3 U34 ( .I(n214), .O(n605) );
  XNR2P U35 ( .I1(n1507), .I2(n1789), .O(n474) );
  XOR2P U36 ( .I1(n2173), .I2(n2124), .O(n471) );
  XOR2P U37 ( .I1(n2254), .I2(n2255), .O(n357) );
  INV3 U38 ( .I(n894), .O(n334) );
  XOR2P U39 ( .I1(n1383), .I2(n1384), .O(n135) );
  INV3 U40 ( .I(n38), .O(n46) );
  OR3B2 U41 ( .I1(n532), .B1(n40), .B2(n1550), .O(n1549) );
  INV2 U42 ( .I(n425), .O(n402) );
  INV2 U43 ( .I(n456), .O(n434) );
  INV2 U44 ( .I(n895), .O(n2008) );
  BUF1 U45 ( .I(n2515), .O(n2507) );
  AOI13HS U46 ( .B1(n474), .B2(n1245), .B3(n471), .A1(n1246), .O(n1244) );
  AOI112P U47 ( .C1(n1541), .C2(n2395), .A1(n1542), .B1(n1543), .O(n1540) );
  XOR2P U48 ( .I1(n1738), .I2(din[26]), .O(n675) );
  NR2T U49 ( .I1(n40), .I2(n539), .O(n1081) );
  XNR2P U50 ( .I1(din[16]), .I2(n1739), .O(n40) );
  AOI13HS U51 ( .B1(n2148), .B2(n474), .B3(n932), .A1(n2149), .O(n2144) );
  INV1 U52 ( .I(n934), .O(n929) );
  AOI13HS U53 ( .B1(n675), .B2(n1811), .B3(n689), .A1(n1812), .O(n1810) );
  BUF1 U54 ( .I(n111), .O(n2424) );
  BUF1 U55 ( .I(n487), .O(n2317) );
  NR2P U56 ( .I1(n2428), .I2(n2431), .O(n417) );
  NR2P U57 ( .I1(n2359), .I2(n2363), .O(n685) );
  INV2 U58 ( .I(n2314), .O(n368) );
  NR2P U59 ( .I1(n2378), .I2(n958), .O(n71) );
  ND2 U60 ( .I1(n548), .I2(n1110), .O(n560) );
  ND2 U61 ( .I1(n2205), .I2(n2280), .O(n1190) );
  BUF1 U62 ( .I(n264), .O(n2390) );
  BUF1 U63 ( .I(n164), .O(n2417) );
  NR2P U64 ( .I1(n582), .I2(n1016), .O(n198) );
  ND3 U65 ( .I1(n361), .I2(n632), .I3(n629), .O(n355) );
  ND2 U66 ( .I1(n1618), .I2(n819), .O(n245) );
  BUF1 U67 ( .I(n480), .O(n2320) );
  BUF1 U68 ( .I(n508), .O(n2330) );
  XNR2 U69 ( .I1(n2181), .I2(n368), .O(n635) );
  BUF1 U70 ( .I(n480), .O(n2321) );
  AOI13HS U71 ( .B1(n307), .B2(n313), .B3(n314), .A1(n315), .O(n296) );
  ND3 U72 ( .I1(n870), .I2(n2340), .I3(n1295), .O(n293) );
  NR2 U73 ( .I1(n451), .I2(n2418), .O(n450) );
  BUF1 U74 ( .I(n427), .O(n2420) );
  OR3 U75 ( .I1(n82), .I2(n1), .I3(n2), .O(n81) );
  OR2 U76 ( .I1(n106), .I2(n107), .O(n1) );
  AO112 U77 ( .C1(n2354), .C2(n86), .A1(n87), .B1(n88), .O(n2) );
  OR3 U78 ( .I1(n55), .I2(n56), .I3(n57), .O(n54) );
  OR2 U79 ( .I1(n79), .I2(n80), .O(n56) );
  AO112 U80 ( .C1(n58), .C2(n2367), .A1(n60), .B1(n61), .O(n57) );
  NR2P U81 ( .I1(n2200), .I2(n2205), .O(n638) );
  NR2P U82 ( .I1(n590), .I2(n1859), .O(n196) );
  NR2P U83 ( .I1(n257), .I2(n814), .O(n1614) );
  NR2P U84 ( .I1(n2415), .I2(n2408), .O(n159) );
  NR2P U85 ( .I1(n2283), .I2(n1740), .O(n1211) );
  NR2P U86 ( .I1(n674), .I2(n101), .O(n989) );
  NR2P U87 ( .I1(n709), .I2(n2378), .O(n957) );
  INV2 U88 ( .I(n275), .O(n285) );
  INV2 U89 ( .I(n247), .O(n257) );
  NR2P U90 ( .I1(n361), .I2(n627), .O(n2205) );
  NR2P U91 ( .I1(n590), .I2(n1029), .O(n1853) );
  INV2 U92 ( .I(n590), .O(n1016) );
  NR2P U93 ( .I1(n2403), .I2(n147), .O(n451) );
  INV2 U94 ( .I(n814), .O(n801) );
  INV2 U95 ( .I(n2354), .O(n689) );
  NR2P U96 ( .I1(n101), .I2(n990), .O(n98) );
  INV2 U97 ( .I(n674), .O(n990) );
  NR2P U98 ( .I1(n382), .I2(n648), .O(n2281) );
  NR2P U99 ( .I1(n285), .I2(n824), .O(n1673) );
  ND3 U100 ( .I1(n1867), .I2(n1868), .I3(n1869), .O(n180) );
  INV2 U101 ( .I(n2404), .O(n158) );
  BUF1 U102 ( .I(n427), .O(n2419) );
  BUF1 U103 ( .I(n486), .O(n2319) );
  ND2 U104 ( .I1(n1321), .I2(n2331), .O(n2019) );
  ND3 U105 ( .I1(n1359), .I2(n1360), .I3(n1361), .O(n751) );
  AOI13HS U106 ( .B1(n2430), .B2(n130), .B3(n757), .A1(n1362), .O(n1361) );
  ND2 U107 ( .I1(n1295), .I2(n1294), .O(n1974) );
  BUF1 U108 ( .I(n427), .O(n2421) );
  ND3 U109 ( .I1(n1156), .I2(n1157), .I3(n1158), .O(n827) );
  ND3 U110 ( .I1(n1129), .I2(n1130), .I3(n1131), .O(n804) );
  XNR2 U111 ( .I1(n275), .I2(n2389), .O(n1169) );
  XNR2 U112 ( .I1(n247), .I2(n236), .O(n1142) );
  ND3 U113 ( .I1(n2385), .I2(n2387), .I3(n2390), .O(n1672) );
  OAI12 U114 ( .B1(n1016), .B2(n1859), .A1(n1025), .O(n193) );
  BUF1 U115 ( .I(n123), .O(n2432) );
  ND2 U116 ( .I1(n129), .I2(n410), .O(n1358) );
  ND3 U117 ( .I1(n1920), .I2(n1921), .I3(n1922), .O(n208) );
  OAI112S U118 ( .C1(n993), .C2(n690), .A1(n994), .B1(n995), .O(n978) );
  MOAI1 U119 ( .A1(n303), .A2(n855), .B1(n309), .B2(n1295), .O(n1305) );
  NR2P U120 ( .I1(n2324), .I2(n512), .O(n914) );
  NR2P U121 ( .I1(n2372), .I2(n62), .O(n718) );
  NR2P U122 ( .I1(n2365), .I2(n2370), .O(n948) );
  NR2P U123 ( .I1(n468), .I2(n489), .O(n934) );
  NR2P U124 ( .I1(n2353), .I2(n2358), .O(n980) );
  NR2P U125 ( .I1(n551), .I2(n22), .O(n1105) );
  INV2 U126 ( .I(n484), .O(n489) );
  INV2 U127 ( .I(n366), .O(n359) );
  INV2 U128 ( .I(n2367), .O(n722) );
  INV2 U129 ( .I(n709), .O(n958) );
  INV2 U130 ( .I(n282), .O(n840) );
  ND3 U131 ( .I1(n135), .I2(n736), .I3(n737), .O(n128) );
  ND2 U132 ( .I1(n101), .I2(n2355), .O(n690) );
  ND3 U133 ( .I1(n1169), .I2(n2388), .I3(n1174), .O(n272) );
  ND2 U134 ( .I1(n2378), .I2(n2368), .O(n724) );
  ND3 U135 ( .I1(n1142), .I2(n252), .I3(n1147), .O(n244) );
  ND2 U136 ( .I1(n1688), .I2(n842), .O(n273) );
  BUF1 U137 ( .I(n369), .O(n2280) );
  XNR2 U138 ( .I1(n309), .I2(n2341), .O(n304) );
  XNR2 U139 ( .I1(n380), .I2(n2006), .O(n656) );
  BUF1 U140 ( .I(n369), .O(n2313) );
  NR2 U141 ( .I1(n2409), .I2(n2405), .O(n787) );
  NR2 U142 ( .I1(n1622), .I2(n2391), .O(n1620) );
  AOI13HS U143 ( .B1(n252), .B2(n811), .B3(n1147), .A1(n241), .O(n1622) );
  AOI13HS U144 ( .B1(n254), .B2(n1148), .B3(n809), .A1(n1149), .O(n1136) );
  AOI13HS U145 ( .B1(n2431), .B2(n2427), .B3(n126), .A1(n127), .O(n115) );
  AOI13HS U146 ( .B1(n627), .B2(n628), .B3(n629), .A1(n630), .O(n626) );
  OAI112S U147 ( .C1(n511), .C2(n918), .A1(n512), .B1(n2329), .O(n917) );
  OAI12S U148 ( .B1(n305), .B2(n303), .A1(n864), .O(n858) );
  NR2P U149 ( .I1(n1042), .I2(n605), .O(n226) );
  ND3 U150 ( .I1(n1817), .I2(n2005), .I3(n1213), .O(n2293) );
  ND2 U151 ( .I1(n282), .I2(n2383), .O(n1172) );
  ND2 U152 ( .I1(n254), .I2(n806), .O(n1145) );
  ND3 U153 ( .I1(n897), .I2(n2335), .I3(n1321), .O(n320) );
  NR2 U154 ( .I1(n1082), .I2(n1083), .O(n1079) );
  ND3 U155 ( .I1(n882), .I2(n323), .I3(n2037), .O(n876) );
  NR2 U156 ( .I1(n319), .I2(n334), .O(n2037) );
  ND3 U157 ( .I1(n614), .I2(n603), .I3(n1906), .O(n1049) );
  ND3 U158 ( .I1(n224), .I2(n603), .I3(n610), .O(n608) );
  ND2 U159 ( .I1(n253), .I2(n1627), .O(n802) );
  XNR2 U160 ( .I1(n897), .I2(n2334), .O(n331) );
  AOI13HS U161 ( .B1(n334), .B2(n340), .B3(n341), .A1(n342), .O(n324) );
  AOI13HS U162 ( .B1(n704), .B2(n2374), .B3(n705), .A1(n78), .O(n700) );
  AOI13HS U163 ( .B1(n648), .B2(n649), .B3(n650), .A1(n651), .O(n647) );
  OAI12S U164 ( .B1(n327), .B2(n328), .A1(n319), .O(n326) );
  NR2 U165 ( .I1(n1111), .I2(n1112), .O(n1108) );
  NR2P U166 ( .I1(n1547), .I2(n525), .O(n41) );
  NR2P U167 ( .I1(n1119), .I2(n548), .O(n18) );
  NR2P U168 ( .I1(n2310), .I2(encrypt_shift[3]), .O(n1446) );
  INV2 U169 ( .I(n1912), .O(n1054) );
  ND2 U170 ( .I1(n548), .I2(n1119), .O(n565) );
  BUF1 U171 ( .I(n515), .O(n2323) );
  BUF1 U172 ( .I(n829), .O(n2385) );
  ND3 U173 ( .I1(n116), .I2(n424), .I3(n2430), .O(n1344) );
  BUF1 U174 ( .I(n813), .O(n2392) );
  BUF1 U175 ( .I(n152), .O(n2416) );
  BUF1 U176 ( .I(n813), .O(n2391) );
  BUF1 U177 ( .I(n66), .O(n2373) );
  BUF1 U178 ( .I(n220), .O(n2349) );
  OAI12 U179 ( .B1(n1042), .B2(n1912), .A1(n1051), .O(n221) );
  BUF1 U180 ( .I(n144), .O(n2408) );
  BUF1 U181 ( .I(n144), .O(n2407) );
  AOI13HS U182 ( .B1(n437), .B2(n170), .B3(n438), .A1(n167), .O(n436) );
  OAI12S U183 ( .B1(n2355), .B2(n691), .A1(n690), .O(n1811) );
  OAI12S U184 ( .B1(n2009), .B2(n337), .A1(n2010), .O(n2007) );
  AOI13HS U185 ( .B1(n2336), .B2(n2333), .B3(n332), .A1(n2013), .O(n2009) );
  NR2P U186 ( .I1(n386), .I2(n1802), .O(n1221) );
  NR2P U187 ( .I1(n613), .I2(n1041), .O(n1050) );
  INV2 U188 ( .I(n386), .O(n374) );
  INV2 U189 ( .I(n16), .O(n551) );
  INV2 U190 ( .I(n613), .O(n1042) );
  INV2 U191 ( .I(n1119), .O(n22) );
  NR2P U192 ( .I1(encrypt_shift[2]), .I2(encrypt_shift[3]), .O(n1448) );
  INV2 U193 ( .I(n837), .O(n824) );
  INV2 U194 ( .I(n655), .O(n382) );
  INV2 U195 ( .I(n25), .O(n563) );
  ND3 U196 ( .I1(n1801), .I2(n386), .I3(n653), .O(n2282) );
  ND3 U197 ( .I1(n768), .I2(n167), .I3(n769), .O(n157) );
  NR2 U198 ( .I1(n2418), .I2(n2405), .O(n769) );
  ND3 U199 ( .I1(n877), .I2(n2333), .I3(n334), .O(n2024) );
  BUF1 U200 ( .I(n59), .O(n2367) );
  BUF1 U201 ( .I(n889), .O(n2334) );
  BUF1 U202 ( .I(n496), .O(n2324) );
  BUF1 U203 ( .I(n813), .O(n2393) );
  BUF1 U204 ( .I(n836), .O(n2381) );
  BUF1 U205 ( .I(n280), .O(n2388) );
  BUF1 U206 ( .I(n514), .O(n2327) );
  BUF1 U207 ( .I(n393), .O(n1961) );
  BUF1 U208 ( .I(n280), .O(n2387) );
  BUF1 U209 ( .I(n829), .O(n2384) );
  BUF1 U210 ( .I(n889), .O(n2336) );
  BUF1 U211 ( .I(n514), .O(n2328) );
  BUF1 U212 ( .I(n708), .O(n2376) );
  BUF1 U213 ( .I(n1320), .O(n2332) );
  BUF1 U214 ( .I(n59), .O(n2365) );
  BUF1 U215 ( .I(n377), .O(n1802) );
  BUF1 U216 ( .I(n390), .O(n1740) );
  BUF1 U217 ( .I(n1320), .O(n2331) );
  BUF1 U218 ( .I(n66), .O(n2372) );
  BUF1 U219 ( .I(n280), .O(n2386) );
  BUF1 U220 ( .I(n708), .O(n2375) );
  AOI13HS U221 ( .B1(n2360), .B2(n670), .B3(n671), .A1(n105), .O(n666) );
  BUF1 U222 ( .I(n144), .O(n2406) );
  AOI13HS U223 ( .B1(n449), .B2(n2405), .B3(n1434), .A1(n1435), .O(n1432) );
  BUF1 U224 ( .I(n836), .O(n2380) );
  MOAI1 U225 ( .A1(n330), .A2(n882), .B1(n337), .B2(n1321), .O(n1331) );
  NR2P U226 ( .I1(n167), .I2(n2410), .O(n793) );
  ND3 U227 ( .I1(n138), .I2(n424), .I3(n416), .O(n425) );
  ND3 U228 ( .I1(n1119), .I2(n25), .I3(n21), .O(n1120) );
  BUF1 U229 ( .I(n514), .O(n2326) );
  BUF1 U230 ( .I(n220), .O(n2348) );
  NR2 U231 ( .I1(n2347), .I2(n1912), .O(n1927) );
  BUF1 U232 ( .I(n708), .O(n2377) );
  BUF1 U233 ( .I(n377), .O(n1960) );
  BUF1 U234 ( .I(n1104), .O(n2399) );
  BUF1 U235 ( .I(n66), .O(n2374) );
  BUF1 U236 ( .I(n1104), .O(n2400) );
  BUF1 U237 ( .I(n390), .O(n1800) );
  BUF1 U238 ( .I(n59), .O(n2366) );
  MOAI1P U239 ( .A1(n2522), .A2(n1937), .B1(n1938), .B2(n2526), .O(n214) );
  INV2 U240 ( .I(din[11]), .O(n1388) );
  BUF1 U241 ( .I(n2554), .O(n2552) );
  INV2 U242 ( .I(n928), .O(n491) );
  INV2 U243 ( .I(n410), .O(n742) );
  INV2 U244 ( .I(n736), .O(n409) );
  INV2 U245 ( .I(n1343), .O(n744) );
  INV2 U246 ( .I(n1184), .O(n2190) );
  INV2 U247 ( .I(n1981), .O(n1304) );
  OAI12 U248 ( .B1(n2424), .B2(n2426), .A1(n746), .O(n736) );
  NR2P U249 ( .I1(n146), .I2(n2409), .O(n443) );
  NR2T U250 ( .I1(n937), .I2(n2317), .O(n928) );
  NR3P U251 ( .I1(n761), .I2(n1354), .I3(n760), .O(n1362) );
  NR2P U252 ( .I1(n116), .I2(n2426), .O(n410) );
  BUF2 U253 ( .I(n2096), .O(n2450) );
  BUF2 U254 ( .I(n2096), .O(n2451) );
  BUF2 U255 ( .I(n2096), .O(n2452) );
  INV2 U256 ( .I(n1018), .O(n592) );
  NR2P U257 ( .I1(n713), .I2(n2370), .O(n953) );
  NR2P U258 ( .I1(n130), .I2(n2431), .O(n1343) );
  BUF2 U259 ( .I(n297), .O(n2341) );
  NR2P U260 ( .I1(n680), .I2(n2357), .O(n985) );
  BUF2 U261 ( .I(n297), .O(n2342) );
  BUF2 U262 ( .I(n111), .O(n2425) );
  BUF1 U263 ( .I(n104), .O(n2361) );
  INV2 U264 ( .I(n560), .O(n9) );
  OR2 U265 ( .I1(n592), .I2(n199), .O(n188) );
  INV2 U266 ( .I(n1602), .O(n811) );
  BUF1 U267 ( .I(n104), .O(n2362) );
  INV2 U268 ( .I(n71), .O(n715) );
  NR2P U269 ( .I1(n725), .I2(n2370), .O(n973) );
  NR2P U270 ( .I1(n691), .I2(n2357), .O(n1005) );
  BUF2 U271 ( .I(n2096), .O(n2453) );
  INV2 U272 ( .I(n419), .O(n423) );
  NR2P U273 ( .I1(n682), .I2(n2362), .O(n1798) );
  INV2 U274 ( .I(n1240), .O(n1238) );
  INV2 U275 ( .I(n635), .O(n636) );
  INV2 U276 ( .I(n1295), .O(n302) );
  OA22 U277 ( .A1(n116), .A2(n759), .B1(n760), .B2(n761), .O(n752) );
  NR2 U278 ( .I1(n1240), .I2(n491), .O(n2149) );
  INV2 U279 ( .I(n1425), .O(n788) );
  INV2 U280 ( .I(n417), .O(n761) );
  INV2 U281 ( .I(n481), .O(n938) );
  NR2 U282 ( .I1(n2430), .I2(n742), .O(n1363) );
  NR2 U283 ( .I1(n71), .I2(n72), .O(n70) );
  INV2 U284 ( .I(n1412), .O(n776) );
  INV2 U285 ( .I(n1741), .O(n961) );
  INV2 U286 ( .I(n685), .O(n996) );
  INV2 U287 ( .I(n1207), .O(n2267) );
  INV2 U288 ( .I(n1803), .O(n993) );
  NR2 U289 ( .I1(n2214), .I2(n630), .O(n2213) );
  INV2 U290 ( .I(n355), .O(n2214) );
  INV2 U291 ( .I(n1289), .O(n1975) );
  INV2 U292 ( .I(n407), .O(n1354) );
  ND2 U293 ( .I1(n2320), .I2(n481), .O(n479) );
  INV2 U294 ( .I(n449), .O(n792) );
  INV2 U295 ( .I(n241), .O(n235) );
  INV2 U296 ( .I(n1188), .O(n2195) );
  INV2 U297 ( .I(n124), .O(n415) );
  OAI12S U298 ( .B1(n312), .B2(n1979), .A1(n849), .O(n1971) );
  NR2P U299 ( .I1(n2431), .I2(n2426), .O(n416) );
  ND2 U300 ( .I1(n1674), .I2(n2390), .O(n1160) );
  OA13 U301 ( .B1(n423), .B2(n2427), .B3(n761), .A1(n405), .O(n1364) );
  INV2 U302 ( .I(n768), .O(n441) );
  INV2 U303 ( .I(n711), .O(n965) );
  NR2 U304 ( .I1(n2337), .I2(n2344), .O(n1300) );
  INV2 U305 ( .I(n629), .O(n1201) );
  ND2 U306 ( .I1(n188), .I2(n1023), .O(n1022) );
  INV2 U307 ( .I(n1276), .O(n907) );
  INV2 U308 ( .I(n170), .O(n166) );
  INV2 U309 ( .I(n269), .O(n263) );
  INV2 U310 ( .I(n293), .O(n1284) );
  INV2 U311 ( .I(n2533), .O(n2521) );
  INV2 U312 ( .I(n2532), .O(n2518) );
  INV2 U313 ( .I(n2532), .O(n2519) );
  INV2 U314 ( .I(n2531), .O(n2517) );
  INV2 U315 ( .I(n2534), .O(n2526) );
  INV2 U316 ( .I(n2531), .O(n2528) );
  INV2 U317 ( .I(n2532), .O(n2529) );
  INV2 U318 ( .I(n2532), .O(n2520) );
  INV2 U319 ( .I(n2533), .O(n2522) );
  INV2 U320 ( .I(n2533), .O(n2523) );
  INV2 U321 ( .I(n2533), .O(n2524) );
  INV2 U322 ( .I(n2533), .O(n2525) );
  INV2 U323 ( .I(n2534), .O(n2527) );
  NR3P U324 ( .I1(n852), .I2(n853), .I3(n854), .O(n295) );
  AO13 U325 ( .B1(n2341), .B2(n855), .B3(n856), .A1(n857), .O(n854) );
  BUF2 U326 ( .I(n292), .O(n2337) );
  INV2 U327 ( .I(n1307), .O(n308) );
  NR2P U328 ( .I1(n2193), .I2(n352), .O(n1184) );
  ND2 U329 ( .I1(n855), .I2(n2339), .O(n1981) );
  NR2 U330 ( .I1(n290), .I2(n291), .O(n289) );
  OAI112S U331 ( .C1(n296), .C2(n2341), .A1(n298), .B1(n299), .O(n290) );
  OAI112S U332 ( .C1(n2337), .C2(n293), .A1(n294), .B1(n295), .O(n291) );
  OAI12S U333 ( .B1(n300), .B2(n301), .A1(n2337), .O(n299) );
  ND2 U334 ( .I1(n622), .I2(n351), .O(n2189) );
  NR3P U335 ( .I1(n359), .I2(n632), .I3(n2315), .O(n1189) );
  NR3P U336 ( .I1(n996), .I2(n689), .I3(n102), .O(n998) );
  NR3P U337 ( .I1(n811), .I2(n809), .I3(n1145), .O(n241) );
  NR3P U338 ( .I1(n534), .I2(n2397), .I3(n36), .O(n35) );
  NR3P U339 ( .I1(n558), .I2(n2402), .I3(n13), .O(n12) );
  NR2T U340 ( .I1(n187), .I2(n176), .O(n587) );
  INV3 U341 ( .I(n2352), .O(n1028) );
  INV3 U342 ( .I(n2181), .O(n352) );
  NR2T U343 ( .I1(n307), .I2(n2343), .O(n1295) );
  OAI112 U344 ( .C1(n2413), .C2(n1415), .A1(n1416), .B1(n780), .O(n168) );
  OR2B1 U345 ( .I1(n1413), .B1(n1422), .O(n1416) );
  AOI13HS U346 ( .B1(n439), .B2(n2412), .B3(n1423), .A1(n1424), .O(n1415) );
  MOAI1 U347 ( .A1(n455), .A2(n2410), .B1(n147), .B2(n1423), .O(n1422) );
  INV2 U348 ( .I(n2420), .O(n130) );
  ND3P U349 ( .I1(n473), .I2(n483), .I3(n489), .O(n1240) );
  ND3P U350 ( .I1(n1016), .I2(n582), .I3(n589), .O(n183) );
  NR2T U351 ( .I1(n1016), .I2(n1029), .O(n1018) );
  OAI12 U352 ( .B1(n2317), .B2(n2319), .A1(n490), .O(n481) );
  INV3 U353 ( .I(n2428), .O(n116) );
  OAI12S U354 ( .B1(n1251), .B2(n2320), .A1(n927), .O(n1250) );
  AOI13HS U355 ( .B1(n483), .B2(n489), .B3(n938), .A1(n1252), .O(n1251) );
  NR2 U356 ( .I1(n483), .I2(n490), .O(n1252) );
  NR2P U357 ( .I1(n870), .I2(n305), .O(n1306) );
  INV3 U358 ( .I(n2411), .O(n146) );
  NR2T U359 ( .I1(n2411), .I2(n2413), .O(n449) );
  AOI13HS U360 ( .B1(n2340), .B2(n869), .B3(n870), .A1(n871), .O(n866) );
  NR2P U361 ( .I1(n491), .I2(n473), .O(n1236) );
  INV2 U362 ( .I(n2319), .O(n937) );
  BUF2 U363 ( .I(n120), .O(n2430) );
  NR2P U364 ( .I1(n2318), .I2(n489), .O(n1249) );
  ND2P U365 ( .I1(n2343), .I2(n307), .O(n303) );
  BUF2 U366 ( .I(n125), .O(n2427) );
  BUF2 U367 ( .I(n120), .O(n2431) );
  OA112 U368 ( .C1(n811), .C2(n1133), .A1(n1612), .B1(n1613), .O(n1127) );
  ND3 U369 ( .I1(n243), .I2(n819), .I3(n1135), .O(n1612) );
  AOI13HS U370 ( .B1(n817), .B2(n1614), .B3(n818), .A1(n1615), .O(n1613) );
  NR3P U371 ( .I1(n1608), .I2(n817), .I3(n246), .O(n1615) );
  BUF2 U372 ( .I(n153), .O(n2409) );
  BUF2 U373 ( .I(n125), .O(n2426) );
  NR2P U374 ( .I1(n257), .I2(n801), .O(n1602) );
  BUF2 U375 ( .I(n73), .O(n2370) );
  OAI112 U376 ( .C1(n2150), .C2(n2151), .A1(n2152), .B1(n2153), .O(n1231) );
  INV2 U377 ( .I(n2147), .O(n2150) );
  ND3 U378 ( .I1(n473), .I2(n1237), .I3(n928), .O(n2152) );
  AOI13HS U379 ( .B1(n2321), .B2(n1236), .B3(n934), .A1(n2154), .O(n2153) );
  XNR2 U380 ( .I1(n2410), .I2(n2412), .O(n1419) );
  NR2P U381 ( .I1(n2417), .I2(n147), .O(n439) );
  BUF2 U382 ( .I(n153), .O(n2410) );
  BUF2 U383 ( .I(n292), .O(n2338) );
  ND3 U384 ( .I1(n990), .I2(n2358), .I3(n673), .O(n995) );
  ND3 U385 ( .I1(n937), .I2(n932), .I3(n2163), .O(n1242) );
  NR2 U386 ( .I1(n2320), .I2(n473), .O(n2163) );
  OAI112 U387 ( .C1(n200), .C2(n1861), .A1(n1862), .B1(n1863), .O(n573) );
  ND3 U388 ( .I1(n587), .I2(n1018), .I3(n1866), .O(n1862) );
  OA22 U389 ( .A1(n1864), .A2(n1015), .B1(n1017), .B2(n1019), .O(n1863) );
  ND3 U390 ( .I1(n582), .I2(n197), .I3(n1024), .O(n577) );
  INV3 U391 ( .I(n2490), .O(n2489) );
  OAI112S U392 ( .C1(n483), .C2(n937), .A1(n489), .B1(n2321), .O(n936) );
  BUF2 U393 ( .I(n100), .O(n2357) );
  OA222 U394 ( .A1(n2209), .A2(n2199), .B1(n2206), .B2(n2210), .C1(n2195), 
        .C2(n2193), .O(n622) );
  OA22 U395 ( .A1(n370), .A2(n2315), .B1(n368), .B2(n637), .O(n2210) );
  INV2 U396 ( .I(n989), .O(n691) );
  INV2 U397 ( .I(n957), .O(n725) );
  NR2P U398 ( .I1(n2421), .I2(n2424), .O(n419) );
  BUF2 U399 ( .I(n100), .O(n2358) );
  NR2P U400 ( .I1(n62), .I2(n77), .O(n1741) );
  ND2P U401 ( .I1(n187), .I2(n1028), .O(n1017) );
  OAI112 U402 ( .C1(n783), .C2(n784), .A1(n785), .B1(n786), .O(n460) );
  INV2 U403 ( .I(n789), .O(n784) );
  ND3 U404 ( .I1(n449), .I2(n159), .I3(n787), .O(n786) );
  OA22 U405 ( .A1(n146), .A2(n790), .B1(n791), .B2(n792), .O(n783) );
  BUF2 U406 ( .I(n553), .O(n2401) );
  BUF2 U407 ( .I(n2092), .O(n2458) );
  ND2P U408 ( .I1(n2316), .I2(n2319), .O(n490) );
  NR2P U409 ( .I1(n2027), .I2(n323), .O(n1330) );
  ND2P U410 ( .I1(n582), .I2(n2352), .O(n199) );
  ND3 U411 ( .I1(n489), .I2(n2164), .I3(n928), .O(n930) );
  BUF2 U412 ( .I(n1375), .O(n2496) );
  BUF2 U413 ( .I(n2090), .O(n2462) );
  BUF2 U414 ( .I(n2094), .O(n2454) );
  ND3 U415 ( .I1(n1028), .I2(n582), .I3(n194), .O(n1861) );
  BUF2 U416 ( .I(n2092), .O(n2459) );
  NR2P U417 ( .I1(n2361), .I2(n2363), .O(n1803) );
  INV2 U418 ( .I(n1095), .O(n558) );
  INV2 U419 ( .I(n1066), .O(n534) );
  BUF2 U420 ( .I(n2094), .O(n2455) );
  BUF2 U421 ( .I(n2092), .O(n2460) );
  BUF2 U422 ( .I(n2090), .O(n2463) );
  BUF2 U423 ( .I(n2094), .O(n2456) );
  BUF2 U424 ( .I(n2090), .O(n2464) );
  BUF2 U425 ( .I(n1377), .O(n2494) );
  INV2 U426 ( .I(n1044), .O(n615) );
  BUF2 U427 ( .I(n487), .O(n2316) );
  AN2B1 U428 ( .I1(n2281), .B1(n380), .O(n1214) );
  NR2P U429 ( .I1(n158), .I2(n2413), .O(n1412) );
  NR2P U430 ( .I1(n2207), .I2(n2181), .O(n1188) );
  OAI12 U431 ( .B1(n62), .B2(n971), .A1(n703), .O(n76) );
  AOI12S U432 ( .B1(n706), .B2(n2378), .A1(n973), .O(n971) );
  NR2P U433 ( .I1(n2432), .I2(n2424), .O(n407) );
  INV2 U434 ( .I(n314), .O(n1290) );
  ND2P U435 ( .I1(n77), .I2(n722), .O(n713) );
  BUF1 U436 ( .I(n529), .O(n2396) );
  AO222 U437 ( .A1(n1184), .A2(n1185), .B1(n1186), .B2(n1187), .C1(n1188), 
        .C2(n1189), .O(n621) );
  OAI12S U438 ( .B1(n2280), .B2(n637), .A1(n1190), .O(n1187) );
  MOAI1P U439 ( .A1(n592), .A2(n2352), .B1(n193), .B2(n2352), .O(n189) );
  MOAI1P U440 ( .A1(n1972), .A2(n2342), .B1(n1306), .B2(n1973), .O(n852) );
  OA22 U441 ( .A1(n1292), .A2(n1974), .B1(n1290), .B2(n1976), .O(n1972) );
  OAI12S U442 ( .B1(n2340), .B2(n1974), .A1(n1975), .O(n1973) );
  INV2 U443 ( .I(n1614), .O(n238) );
  BUF2 U444 ( .I(n311), .O(n2343) );
  ND2P U445 ( .I1(n689), .I2(n2362), .O(n680) );
  NR2P U446 ( .I1(n429), .I2(n751), .O(n132) );
  BUF2 U447 ( .I(n529), .O(n2397) );
  ND2 U448 ( .I1(n1237), .I2(n937), .O(n475) );
  ND2 U449 ( .I1(n1262), .I2(n918), .O(n503) );
  NR2P U450 ( .I1(n180), .I2(n573), .O(n1011) );
  NR2P U451 ( .I1(n208), .I2(n596), .O(n1036) );
  INV2 U452 ( .I(n1673), .O(n834) );
  AO112 U453 ( .C1(n948), .C2(n707), .A1(n949), .B1(n719), .O(n80) );
  AO112 U454 ( .C1(n980), .C2(n673), .A1(n981), .B1(n686), .O(n107) );
  OAI112S U455 ( .C1(n199), .C2(n1025), .A1(n1026), .B1(n1027), .O(n1020) );
  ND3 U456 ( .I1(n582), .I2(n193), .I3(n176), .O(n1026) );
  AOI13HS U457 ( .B1(n1028), .B2(n1029), .B3(n1030), .A1(n1031), .O(n1027) );
  AOI112P U458 ( .C1(n592), .C2(n1032), .A1(n582), .B1(n176), .O(n1031) );
  NR2P U459 ( .I1(n490), .I2(n473), .O(n2143) );
  OAI112S U460 ( .C1(n1017), .C2(n1856), .A1(n1857), .B1(n1858), .O(n1855) );
  INV2 U461 ( .I(n1030), .O(n1856) );
  ND3 U462 ( .I1(n2352), .I2(n592), .I3(n194), .O(n1858) );
  ND3 U463 ( .I1(n1028), .I2(n193), .I3(n587), .O(n1857) );
  INV2 U464 ( .I(n196), .O(n200) );
  INV2 U465 ( .I(n98), .O(n682) );
  OAI12S U466 ( .B1(n2371), .B2(n2379), .A1(n75), .O(n69) );
  ND2P U467 ( .I1(n1306), .I2(n2339), .O(n1979) );
  INV2 U468 ( .I(n268), .O(n1674) );
  ND2P U469 ( .I1(n2311), .I2(n2312), .O(n2096) );
  INV2 U470 ( .I(n240), .O(n1603) );
  NR2P U471 ( .I1(n2270), .I2(n380), .O(n1207) );
  OAI12S U472 ( .B1(n532), .B2(n534), .A1(n535), .O(n530) );
  NR2P U473 ( .I1(n804), .I2(n1128), .O(n250) );
  OAI12S U474 ( .B1(n556), .B2(n558), .A1(n559), .O(n554) );
  INV2 U475 ( .I(n819), .O(n1598) );
  NR2P U476 ( .I1(n827), .I2(n1155), .O(n278) );
  ND2 U477 ( .I1(n2205), .I2(n352), .O(n2199) );
  BUF2 U478 ( .I(n2092), .O(n2461) );
  INV2 U479 ( .I(n1161), .O(n274) );
  BUF2 U480 ( .I(n2094), .O(n2457) );
  BUF2 U481 ( .I(n2090), .O(n2465) );
  NR2P U482 ( .I1(n1976), .I2(n2339), .O(n1289) );
  INV2 U483 ( .I(n932), .O(n478) );
  ND2 U484 ( .I1(n1865), .I2(n176), .O(n1015) );
  ND3 U485 ( .I1(n2427), .I2(n2429), .I3(n1343), .O(n1345) );
  ND2 U486 ( .I1(n818), .I2(n819), .O(n255) );
  NR2P U487 ( .I1(n227), .I2(n204), .O(n1924) );
  NR2P U488 ( .I1(n715), .I2(n77), .O(n1736) );
  NR2P U489 ( .I1(n199), .I2(n176), .O(n1871) );
  ND2 U490 ( .I1(n1134), .I2(n236), .O(n239) );
  ND3 U491 ( .I1(n2313), .I2(n2315), .I3(n638), .O(n367) );
  ND2 U492 ( .I1(n1423), .I2(n2413), .O(n790) );
  NR2P U493 ( .I1(n75), .I2(n2370), .O(n72) );
  INV2 U494 ( .I(n1356), .O(n760) );
  NR2P U495 ( .I1(n621), .I2(n1183), .O(n350) );
  ND2 U496 ( .I1(n1356), .I2(n2430), .O(n759) );
  INV2 U497 ( .I(n908), .O(n518) );
  INV2 U498 ( .I(n1672), .O(n841) );
  NR2P U499 ( .I1(n102), .I2(n2358), .O(n99) );
  INV2 U500 ( .I(n2209), .O(n1186) );
  ND2 U501 ( .I1(n380), .I2(n2281), .O(n2275) );
  INV2 U502 ( .I(n536), .O(n32) );
  INV2 U503 ( .I(n1301), .O(n1292) );
  OR2 U504 ( .I1(n488), .I2(n483), .O(n927) );
  NR2P U505 ( .I1(n939), .I2(n1231), .O(n466) );
  ND2 U506 ( .I1(n1603), .I2(n236), .O(n1133) );
  ND2 U507 ( .I1(n159), .I2(n443), .O(n1425) );
  INV2 U508 ( .I(n1185), .O(n2207) );
  AN3 U509 ( .I1(n361), .I2(n2313), .I3(n1189), .O(n630) );
  NR2 U510 ( .I1(n62), .I2(n958), .O(n954) );
  INV2 U511 ( .I(n1799), .O(n992) );
  INV2 U512 ( .I(n248), .O(n1618) );
  INV2 U513 ( .I(n276), .O(n1688) );
  OR3B2 U514 ( .I1(n857), .B1(n294), .B2(n851), .O(n1285) );
  INV2 U515 ( .I(n1737), .O(n960) );
  INV2 U516 ( .I(n1853), .O(n1025) );
  NR2 U517 ( .I1(n2316), .I2(n2151), .O(n2158) );
  INV2 U518 ( .I(n815), .O(n1135) );
  ND3 U519 ( .I1(n183), .I2(n188), .I3(n1860), .O(n1854) );
  ND3 U520 ( .I1(n187), .I2(n197), .I3(n198), .O(n1860) );
  NR2 U521 ( .I1(n187), .I2(n196), .O(n195) );
  NR3P U522 ( .I1(n232), .I2(n233), .I3(n234), .O(n231) );
  OAI112S U523 ( .C1(n242), .C2(n243), .A1(n244), .B1(n245), .O(n233) );
  ND3 U524 ( .I1(n249), .I2(n250), .I3(n251), .O(n232) );
  NR3P U525 ( .I1(n260), .I2(n261), .I3(n262), .O(n259) );
  OAI112S U526 ( .C1(n270), .C2(n271), .A1(n272), .B1(n273), .O(n261) );
  ND3 U527 ( .I1(n277), .I2(n278), .I3(n279), .O(n260) );
  OA112 U528 ( .C1(n1292), .C2(n1975), .A1(n1977), .B1(n1978), .O(n851) );
  ND3 U529 ( .I1(n2342), .I2(n1306), .I3(n856), .O(n1978) );
  AO12 U530 ( .B1(n1291), .B2(n1976), .A1(n1979), .O(n1977) );
  NR2 U531 ( .I1(n990), .I2(n2364), .O(n986) );
  NR2P U532 ( .I1(n642), .I2(n1206), .O(n396) );
  INV2 U533 ( .I(n1265), .O(n1263) );
  NR2 U534 ( .I1(n134), .I2(n430), .O(n1339) );
  NR2 U535 ( .I1(n168), .I2(n461), .O(n1408) );
  NR2 U536 ( .I1(n750), .I2(n430), .O(n749) );
  INV2 U537 ( .I(n132), .O(n750) );
  NR2 U538 ( .I1(n169), .I2(n461), .O(n781) );
  INV2 U539 ( .I(n1291), .O(n1288) );
  INV2 U540 ( .I(n2151), .O(n2142) );
  NR2 U541 ( .I1(n1265), .I2(n518), .O(n2068) );
  INV2 U542 ( .I(n1134), .O(n246) );
  INV2 U543 ( .I(n1358), .O(n757) );
  OR2 U544 ( .I1(n542), .I2(n1065), .O(n50) );
  OR2 U545 ( .I1(n566), .I2(n1094), .O(n26) );
  INV2 U546 ( .I(n1321), .O(n329) );
  ND2 U547 ( .I1(n1127), .I2(n249), .O(n803) );
  ND2 U548 ( .I1(n1154), .I2(n277), .O(n826) );
  INV2 U549 ( .I(n2216), .O(n362) );
  INV2 U550 ( .I(n1543), .O(n535) );
  INV2 U551 ( .I(n1477), .O(n559) );
  NR2 U552 ( .I1(n532), .I2(n533), .O(n531) );
  OR2B1 U553 ( .I1(n460), .B1(n782), .O(n169) );
  ND2 U554 ( .I1(n1197), .I2(n368), .O(n2196) );
  NR2 U555 ( .I1(n174), .I2(n175), .O(n173) );
  OAI112S U556 ( .C1(n181), .C2(n182), .A1(n183), .B1(n184), .O(n174) );
  OAI112S U557 ( .C1(n176), .C2(n177), .A1(n178), .B1(n179), .O(n175) );
  INV2 U558 ( .I(n194), .O(n182) );
  INV2 U559 ( .I(n509), .O(n919) );
  NR2 U560 ( .I1(n571), .I2(n572), .O(n570) );
  ND3 U561 ( .I1(n585), .I2(n177), .I3(n586), .O(n571) );
  OR3B2 U562 ( .I1(n573), .B1(n178), .B2(n574), .O(n572) );
  AOI13HS U563 ( .B1(n582), .B2(n189), .B3(n587), .A1(n588), .O(n586) );
  NR2 U564 ( .I1(n744), .I2(n2422), .O(n1351) );
  NR2 U565 ( .I1(n2426), .I2(n2419), .O(n756) );
  NR2 U566 ( .I1(n1282), .I2(n1283), .O(n1281) );
  OAI112S U567 ( .C1(n1296), .C2(n2339), .A1(n1297), .B1(n1298), .O(n1282) );
  AO112 U568 ( .C1(n305), .C2(n1284), .A1(n853), .B1(n1285), .O(n1283) );
  AOI13HS U569 ( .B1(n865), .B2(n1299), .B3(n1300), .A1(n301), .O(n1298) );
  INV2 U570 ( .I(n1558), .O(n1067) );
  AN2 U571 ( .I1(n583), .I2(n584), .O(n178) );
  NR2 U572 ( .I1(n98), .I2(n99), .O(n97) );
  INV2 U573 ( .I(n1367), .O(n746) );
  NR2 U574 ( .I1(n2419), .I2(n1358), .O(n1357) );
  ND2 U575 ( .I1(n643), .I2(n395), .O(n2266) );
  INV2 U576 ( .I(n683), .O(n979) );
  INV2 U577 ( .I(n716), .O(n947) );
  AN2 U578 ( .I1(n672), .I2(n673), .O(n105) );
  INV2 U579 ( .I(n1232), .O(n923) );
  INV2 U580 ( .I(n1257), .O(n903) );
  NR2 U581 ( .I1(n2199), .I2(n2314), .O(n2202) );
  AO222 U582 ( .A1(n1103), .A2(n1490), .B1(n1491), .B2(n1107), .C1(n1096), 
        .C2(n1110), .O(n1094) );
  OAI12S U583 ( .B1(n2402), .B2(n557), .A1(n14), .O(n1490) );
  NR2 U584 ( .I1(n558), .I2(n1493), .O(n1491) );
  AN3 U585 ( .I1(n449), .I2(n439), .I3(n1423), .O(n1429) );
  AN3 U586 ( .I1(n718), .I2(n956), .I3(n957), .O(n955) );
  AN3 U587 ( .I1(n685), .I2(n988), .I3(n989), .O(n987) );
  INV2 U588 ( .I(n180), .O(n179) );
  INV2 U589 ( .I(n208), .O(n207) );
  INV2 U590 ( .I(n134), .O(n133) );
  INV2 U591 ( .I(n1315), .O(n2020) );
  INV2 U592 ( .I(n751), .O(n1338) );
  ND2 U593 ( .I1(n2330), .I2(n509), .O(n507) );
  INV2 U594 ( .I(n2340), .O(n297) );
  INV2 U595 ( .I(n2359), .O(n104) );
  ND2 U596 ( .I1(n840), .I2(n1673), .O(n1677) );
  INV2 U597 ( .I(n2422), .O(n111) );
  INV2 U598 ( .I(n1554), .O(n1074) );
  INV2 U599 ( .I(n1488), .O(n1103) );
  OR2 U600 ( .I1(n430), .I2(n134), .O(n428) );
  OR2 U601 ( .I1(n461), .I2(n168), .O(n459) );
  XNR2 U602 ( .I1(n2419), .I2(n2429), .O(n138) );
  NR3P U603 ( .I1(n964), .I2(n722), .I3(n75), .O(n966) );
  ND3P U604 ( .I1(n116), .I2(n2421), .I3(n2433), .O(n124) );
  NR3P U605 ( .I1(n834), .I2(n831), .I3(n1172), .O(n269) );
  AOI112P U606 ( .C1(n302), .C2(n303), .A1(n304), .B1(n305), .O(n300) );
  ND3P U607 ( .I1(n187), .I2(n1018), .I3(n1866), .O(n177) );
  OAI12 U608 ( .B1(n147), .B2(n2409), .A1(n778), .O(n768) );
  NR2T U609 ( .I1(n2181), .I2(n359), .O(n629) );
  ND3P U610 ( .I1(n2379), .I2(n956), .I3(n1741), .O(n711) );
  INV3 U611 ( .I(n2490), .O(n2487) );
  INV3 U612 ( .I(n2485), .O(n2482) );
  AOI112P U613 ( .C1(n2401), .C2(n9), .A1(n1477), .B1(n1478), .O(n1476) );
  NR2 U614 ( .I1(n548), .I2(n14), .O(n1478) );
  XNR2 U615 ( .I1(n729), .I2(n2378), .O(n1754) );
  INV3 U616 ( .I(n2475), .O(n2471) );
  INV3 U617 ( .I(n2490), .O(n2488) );
  ND3P U618 ( .I1(n116), .I2(n2419), .I3(n762), .O(n137) );
  BUF2 U619 ( .I(n1375), .O(n2495) );
  INV3 U620 ( .I(n2485), .O(n2483) );
  INV3 U621 ( .I(n2470), .O(n2466) );
  BUF2 U622 ( .I(n73), .O(n2371) );
  ND3 U623 ( .I1(n958), .I2(n2371), .I3(n707), .O(n963) );
  INV3 U624 ( .I(n2474), .O(n2472) );
  BUF2 U625 ( .I(n1377), .O(n2492) );
  INV3 U626 ( .I(n2469), .O(n2467) );
  INV3 U627 ( .I(n2485), .O(n2484) );
  ND3 U628 ( .I1(n1028), .I2(n591), .I3(n1853), .O(n1023) );
  INV2 U629 ( .I(n442), .O(n154) );
  BUF2 U630 ( .I(n1442), .O(n2479) );
  ND3 U631 ( .I1(n1028), .I2(n196), .I3(n587), .O(n585) );
  BUF2 U632 ( .I(n553), .O(n2402) );
  BUF2 U633 ( .I(n1377), .O(n2493) );
  BUF2 U634 ( .I(n1444), .O(n2476) );
  ND3 U635 ( .I1(n2433), .I2(n762), .I3(n763), .O(n121) );
  NR2 U636 ( .I1(n2420), .I2(n2428), .O(n763) );
  ND3 U637 ( .I1(n443), .I2(n147), .I3(n444), .O(n170) );
  NR2 U638 ( .I1(n158), .I2(n2417), .O(n444) );
  OAI12 U639 ( .B1(n990), .B2(n677), .A1(n676), .O(n82) );
  BUF2 U640 ( .I(n1442), .O(n2480) );
  BUF2 U641 ( .I(n1375), .O(n2497) );
  OAI12 U642 ( .B1(n958), .B2(n711), .A1(n710), .O(n55) );
  BUF2 U643 ( .I(n1444), .O(n2477) );
  INV2 U644 ( .I(n2475), .O(n2473) );
  ND3 U645 ( .I1(n1803), .I2(n988), .I3(n989), .O(n676) );
  ND3 U646 ( .I1(n1741), .I2(n956), .I3(n957), .O(n710) );
  ND3 U647 ( .I1(n2342), .I2(n855), .I3(n1987), .O(n849) );
  NR2 U648 ( .I1(n2337), .I2(n307), .O(n1987) );
  INV2 U649 ( .I(n2470), .O(n2468) );
  BUF1 U650 ( .I(n508), .O(n2329) );
  ND3 U651 ( .I1(n2425), .I2(n410), .I3(n411), .O(n131) );
  NR2 U652 ( .I1(n130), .I2(n2432), .O(n411) );
  ND3 U653 ( .I1(n2338), .I2(n314), .I3(n1295), .O(n868) );
  ND3 U654 ( .I1(n147), .I2(n2412), .I3(n1423), .O(n437) );
  ND3 U655 ( .I1(n138), .I2(n2433), .I3(n139), .O(n136) );
  NR2P U656 ( .I1(n516), .I2(n511), .O(n1276) );
  OAI112S U657 ( .C1(n1144), .C2(n1145), .A1(n1146), .B1(n253), .O(n1143) );
  ND3 U658 ( .I1(n236), .I2(n257), .I3(n1147), .O(n1146) );
  INV2 U659 ( .I(n1142), .O(n1144) );
  OR2 U660 ( .I1(n615), .I2(n227), .O(n216) );
  OAI112S U661 ( .C1(n1171), .C2(n1172), .A1(n1173), .B1(n281), .O(n1170) );
  ND3 U662 ( .I1(n2389), .I2(n285), .I3(n1174), .O(n1173) );
  INV2 U663 ( .I(n1169), .O(n1171) );
  NR2P U664 ( .I1(n582), .I2(n1028), .O(n1866) );
  OAI12S U665 ( .B1(n1614), .B2(n237), .A1(n245), .O(n1619) );
  BUF2 U666 ( .I(n1442), .O(n2481) );
  BUF2 U667 ( .I(n1444), .O(n2478) );
  BUF1 U668 ( .I(n164), .O(n2418) );
  BUF1 U669 ( .I(n264), .O(n2389) );
  MAOI1 U670 ( .A1(n197), .A2(n198), .B1(n199), .B2(n200), .O(n181) );
  BUF1 U671 ( .I(n311), .O(n2344) );
  ND3 U672 ( .I1(n2425), .I2(n2429), .I3(n1356), .O(n405) );
  ND3 U673 ( .I1(n2344), .I2(n1303), .I3(n1304), .O(n1297) );
  NR2P U674 ( .I1(n2413), .I2(n2409), .O(n448) );
  OAI12S U675 ( .B1(n339), .B2(n2025), .A1(n876), .O(n2016) );
  ND3 U676 ( .I1(n2410), .I2(n2412), .I3(n1412), .O(n1414) );
  NR2P U677 ( .I1(n139), .I2(n762), .O(n420) );
  INV2 U678 ( .I(n838), .O(n1162) );
  ND3 U679 ( .I1(n2423), .I2(n741), .I3(n2431), .O(n740) );
  MOAI1 U680 ( .A1(n742), .A2(n130), .B1(n2427), .B2(n415), .O(n741) );
  INV2 U681 ( .I(n1197), .O(n624) );
  INV2 U682 ( .I(n451), .O(n455) );
  INV2 U683 ( .I(n2285), .O(n1209) );
  OR3 U684 ( .I1(n1145), .I2(n238), .I3(n236), .O(n816) );
  OR3 U685 ( .I1(n1172), .I2(n266), .I3(n2389), .O(n839) );
  ND2 U686 ( .I1(n1161), .I2(n2389), .O(n267) );
  INV2 U687 ( .I(n914), .O(n909) );
  INV2 U688 ( .I(n1329), .O(n339) );
  AN3 U689 ( .I1(n159), .I2(n2412), .I3(n162), .O(n457) );
  INV2 U690 ( .I(n1303), .O(n312) );
  INV2 U691 ( .I(n1423), .O(n791) );
  INV2 U692 ( .I(n656), .O(n657) );
  ND3 U693 ( .I1(n445), .I2(n446), .I3(n447), .O(n435) );
  ND3 U694 ( .I1(n2410), .I2(n449), .I3(n450), .O(n446) );
  ND3 U695 ( .I1(n154), .I2(n147), .I3(n448), .O(n447) );
  OR3B2 U696 ( .I1(n452), .B1(n2412), .B2(n454), .O(n445) );
  INV2 U697 ( .I(n1024), .O(n1864) );
  NR2 U698 ( .I1(n556), .I2(n557), .O(n555) );
  INV2 U699 ( .I(n2293), .O(n392) );
  INV2 U700 ( .I(n677), .O(n997) );
  INV2 U701 ( .I(n304), .O(n1299) );
  INV2 U702 ( .I(n331), .O(n1325) );
  NR2 U703 ( .I1(n158), .I2(n159), .O(n155) );
  NR2 U704 ( .I1(n419), .I2(n2433), .O(n418) );
  INV2 U705 ( .I(n1434), .O(n778) );
  AN3 U706 ( .I1(n2344), .I2(n1301), .I3(n1302), .O(n301) );
  NR2 U707 ( .I1(n307), .I2(n2342), .O(n1302) );
  INV2 U708 ( .I(n1492), .O(n1096) );
  INV2 U709 ( .I(n718), .O(n964) );
  ND2 U710 ( .I1(n196), .I2(n192), .O(n1032) );
  AN2 U711 ( .I1(n706), .I2(n707), .O(n78) );
  INV2 U712 ( .I(n650), .O(n1225) );
  ND2 U713 ( .I1(n216), .I2(n1049), .O(n1048) );
  NR2 U714 ( .I1(n2291), .I2(n651), .O(n2290) );
  INV2 U715 ( .I(n379), .O(n2291) );
  INV2 U716 ( .I(n349), .O(n2188) );
  AOI112P U717 ( .C1(n154), .C2(n2414), .A1(n160), .B1(n161), .O(n143) );
  AN3 U718 ( .I1(n162), .I2(n163), .I3(n2417), .O(n161) );
  INV2 U719 ( .I(n165), .O(n160) );
  INV2 U720 ( .I(n526), .O(n1080) );
  INV2 U721 ( .I(n320), .O(n1311) );
  INV2 U722 ( .I(n2508), .O(n2499) );
  INV2 U723 ( .I(n2508), .O(n2500) );
  INV2 U724 ( .I(n2508), .O(n2502) );
  INV2 U725 ( .I(n2508), .O(n2503) );
  INV2 U726 ( .I(n2507), .O(n2501) );
  INV2 U727 ( .I(n2507), .O(n2498) );
  INV2 U728 ( .I(n2508), .O(n2504) );
  BUF1 U729 ( .I(n2538), .O(n2530) );
  BUF2 U730 ( .I(n2537), .O(n2532) );
  BUF2 U731 ( .I(n2537), .O(n2533) );
  BUF2 U732 ( .I(n2536), .O(n2534) );
  BUF1 U733 ( .I(n2538), .O(n2531) );
  BUF1 U734 ( .I(n2536), .O(n2535) );
  MAOI1 U735 ( .A1(n225), .A2(n226), .B1(n227), .B2(n228), .O(n209) );
  INV2 U736 ( .I(n394), .O(n2265) );
  INV2 U737 ( .I(n549), .O(n1109) );
  AOI112P U738 ( .C1(n1186), .C2(n1188), .A1(n1182), .B1(n2197), .O(n351) );
  ND2 U739 ( .I1(n2200), .I2(n2313), .O(n2198) );
  INV3 U740 ( .I(n862), .O(n305) );
  NR2T U741 ( .I1(n309), .I2(n305), .O(n855) );
  ND3P U742 ( .I1(n368), .I2(n357), .I3(n359), .O(n2193) );
  BUF2 U743 ( .I(n2172), .O(n2434) );
  NR2P U744 ( .I1(n850), .I2(n2337), .O(n1307) );
  BUF2 U745 ( .I(n2171), .O(n2440) );
  BUF2 U746 ( .I(n2172), .O(n2436) );
  NR2P U747 ( .I1(n308), .I2(n867), .O(n1983) );
  INV2 U748 ( .I(n1294), .O(n292) );
  BUF2 U749 ( .I(n2171), .O(n2441) );
  BUF2 U750 ( .I(n2172), .O(n2437) );
  AO222 U751 ( .A1(n2342), .A2(n1984), .B1(n1985), .B2(n1304), .C1(n1986), 
        .C2(n1983), .O(n857) );
  NR2 U752 ( .I1(n302), .I2(n1294), .O(n1985) );
  INV2 U753 ( .I(n1979), .O(n1986) );
  MOAI1 U754 ( .A1(n1974), .A2(n1290), .B1(n1301), .B2(n1983), .O(n1984) );
  ND3 U755 ( .I1(n846), .I2(n847), .I3(n848), .O(n845) );
  AOI13HS U756 ( .B1(n309), .B2(n858), .B3(n2338), .A1(n859), .O(n847) );
  OA22 U757 ( .A1(n866), .A2(n867), .B1(n2340), .B2(n868), .O(n846) );
  OA112 U758 ( .C1(n849), .C2(n850), .A1(n851), .B1(n295), .O(n848) );
  ND3 U759 ( .I1(n2185), .I2(n2186), .I3(n2187), .O(n2184) );
  OA22 U760 ( .A1(n1201), .A2(n2216), .B1(n2280), .B2(n353), .O(n2185) );
  OA222 U761 ( .A1(n2211), .A2(n359), .B1(n366), .B2(n2212), .C1(n627), .C2(
        n2213), .O(n2186) );
  AOI112P U762 ( .C1(n2188), .C2(n2314), .A1(n2189), .B1(n1183), .O(n2187) );
  NR3P U763 ( .I1(n483), .I2(n489), .I3(n485), .O(n1237) );
  NR3P U764 ( .I1(n512), .I2(n511), .I3(n2328), .O(n1262) );
  NR3P U765 ( .I1(n809), .I2(n243), .I3(n2392), .O(n818) );
  NR3P U766 ( .I1(n1028), .I2(n582), .I3(n1859), .O(n1865) );
  XNR2 U767 ( .I1(n1859), .I2(n1028), .O(n197) );
  ND3P U768 ( .I1(n563), .I2(n17), .I3(n2401), .O(n14) );
  NR3P U769 ( .I1(n2343), .I2(n2338), .I3(n867), .O(n856) );
  XNR2 U770 ( .I1(n483), .I2(n471), .O(n2164) );
  NR3P U771 ( .I1(n725), .I2(n77), .I3(n2376), .O(n959) );
  AOI112P U772 ( .C1(n1209), .C2(n1211), .A1(n1205), .B1(n2272), .O(n395) );
  ND2 U773 ( .I1(n2276), .I2(n1740), .O(n2274) );
  INV2 U774 ( .I(n2271), .O(n2273) );
  XNR2 U775 ( .I1(n2324), .I2(n500), .O(n2083) );
  INV3 U776 ( .I(n580), .O(n187) );
  INV3 U777 ( .I(n468), .O(n483) );
  ND3P U778 ( .I1(n101), .I2(n674), .I3(n2364), .O(n1799) );
  NR3P U779 ( .I1(n653), .I2(n374), .I3(n2006), .O(n1212) );
  ND3P U780 ( .I1(n2378), .I2(n709), .I3(n62), .O(n1737) );
  NR3P U781 ( .I1(n862), .I2(n308), .I3(n304), .O(n871) );
  INV3 U782 ( .I(n2335), .O(n323) );
  INV3 U783 ( .I(n2375), .O(n62) );
  INV3 U784 ( .I(n2333), .O(n319) );
  INV3 U785 ( .I(n1801), .O(n380) );
  AOI112P U786 ( .C1(n991), .C2(n980), .A1(n88), .B1(n1794), .O(n683) );
  AO13 U787 ( .B1(n2361), .B2(n988), .B3(n992), .A1(n1795), .O(n1794) );
  ND2 U788 ( .I1(n1796), .I2(n1797), .O(n1795) );
  ND3 U789 ( .I1(n2364), .I2(n985), .I3(n1004), .O(n1797) );
  INV3 U790 ( .I(n867), .O(n307) );
  NR2T U791 ( .I1(n801), .I2(n247), .O(n1134) );
  INV3 U792 ( .I(n2407), .O(n147) );
  INV3 U793 ( .I(n2373), .O(n77) );
  INV3 U794 ( .I(n252), .O(n809) );
  NR2T U795 ( .I1(n814), .I2(n247), .O(n819) );
  AOI13HS U796 ( .B1(n2340), .B2(n862), .B3(n2338), .A1(n1970), .O(n1969) );
  NR2 U797 ( .I1(n862), .I2(n2339), .O(n1970) );
  NR2T U798 ( .I1(n2419), .I2(n122), .O(n1356) );
  INV3 U799 ( .I(n806), .O(n243) );
  NR2T U800 ( .I1(n204), .I2(n215), .O(n610) );
  NR2T U801 ( .I1(n334), .I2(n338), .O(n1321) );
  OAI112 U802 ( .C1(n1346), .C2(n2431), .A1(n1347), .B1(n748), .O(n134) );
  ND2 U803 ( .I1(n1352), .I2(n1355), .O(n1347) );
  AOI13HS U804 ( .B1(n407), .B2(n2429), .B3(n1356), .A1(n1357), .O(n1346) );
  MOAI1 U805 ( .A1(n423), .A2(n2427), .B1(n2425), .B2(n1356), .O(n1355) );
  INV3 U806 ( .I(n2345), .O(n204) );
  NR2T U807 ( .I1(n366), .I2(n357), .O(n1197) );
  ND3 U808 ( .I1(n674), .I2(n670), .I3(n688), .O(n95) );
  NR2 U809 ( .I1(n689), .I2(n2361), .O(n688) );
  NR2T U810 ( .I1(n275), .I2(n824), .O(n1161) );
  INV3 U811 ( .I(n2350), .O(n176) );
  INV3 U812 ( .I(n471), .O(n473) );
  OAI12 U813 ( .B1(n513), .B2(n2323), .A1(n517), .O(n509) );
  ND3 U814 ( .I1(n709), .I2(n704), .I3(n721), .O(n68) );
  NR2 U815 ( .I1(n77), .I2(n722), .O(n721) );
  INV3 U816 ( .I(n2386), .O(n831) );
  INV2 U817 ( .I(n17), .O(n1112) );
  INV3 U818 ( .I(n1802), .O(n653) );
  NR2T U819 ( .I1(n17), .I2(n563), .O(n1110) );
  NR2T U820 ( .I1(n2350), .I2(n187), .O(n194) );
  ND3P U821 ( .I1(n483), .I2(n471), .I3(n2159), .O(n2151) );
  NR2 U822 ( .I1(n484), .I2(n2318), .O(n2159) );
  INV3 U823 ( .I(n2349), .O(n603) );
  OR2 U824 ( .I1(n83), .I2(n84), .O(n431) );
  AO112 U825 ( .C1(n457), .C2(n2405), .A1(n459), .B1(n460), .O(n83) );
  AO112 U826 ( .C1(n434), .C2(n2407), .A1(n435), .B1(n436), .O(n84) );
  INV3 U827 ( .I(n2325), .O(n511) );
  INV3 U828 ( .I(n357), .O(n632) );
  INV3 U829 ( .I(n2385), .O(n270) );
  NR2T U830 ( .I1(n2345), .I2(n215), .O(n222) );
  OAI112 U831 ( .C1(n2155), .C2(n2321), .A1(n2156), .B1(n2157), .O(n939) );
  ND3 U832 ( .I1(n2148), .I2(n2147), .I3(n932), .O(n2157) );
  ND3 U833 ( .I1(n2320), .I2(n2316), .I3(n2142), .O(n2156) );
  AOI13HS U834 ( .B1(n468), .B2(n484), .B3(n1236), .A1(n2158), .O(n2155) );
  ND3P U835 ( .I1(n2392), .I2(n254), .I3(n809), .O(n815) );
  ND3P U836 ( .I1(n236), .I2(n254), .I3(n809), .O(n248) );
  INV3 U837 ( .I(n2391), .O(n236) );
  ND3P U838 ( .I1(n500), .I2(n512), .I3(n511), .O(n1265) );
  ND3P U839 ( .I1(n2390), .I2(n282), .I3(n831), .O(n276) );
  INV3 U840 ( .I(n2398), .O(n548) );
  NR2T U841 ( .I1(n1017), .I2(n1859), .O(n589) );
  NR2T U842 ( .I1(n806), .I2(n254), .O(n1147) );
  NR3P U843 ( .I1(n1413), .I2(n147), .I3(n774), .O(n1421) );
  ND3 U844 ( .I1(n366), .I2(n2280), .I3(n632), .O(n2206) );
  ND3 U845 ( .I1(n798), .I2(n799), .I3(n800), .O(n797) );
  OA22 U846 ( .A1(n252), .A2(n816), .B1(n817), .B2(n255), .O(n798) );
  OA222 U847 ( .A1(n805), .A2(n806), .B1(n248), .B2(n807), .C1(n808), .C2(n809), .O(n799) );
  AOI112P U848 ( .C1(n801), .C2(n802), .A1(n803), .B1(n804), .O(n800) );
  ND3 U849 ( .I1(n821), .I2(n822), .I3(n823), .O(n820) );
  OA22 U850 ( .A1(n2388), .A2(n839), .B1(n840), .B2(n283), .O(n821) );
  OA222 U851 ( .A1(n828), .A2(n2384), .B1(n276), .B2(n830), .C1(n831), .C2(
        n832), .O(n822) );
  AOI112P U852 ( .C1(n824), .C2(n825), .A1(n826), .B1(n827), .O(n823) );
  AOI112P U853 ( .C1(n471), .C2(n1247), .A1(n929), .B1(n485), .O(n1246) );
  OAI112S U854 ( .C1(n937), .C2(n478), .A1(n488), .B1(n1248), .O(n1245) );
  ND2 U855 ( .I1(n937), .I2(n2316), .O(n1247) );
  INV2 U856 ( .I(n634), .O(n361) );
  ND3 U857 ( .I1(n484), .I2(n481), .I3(n2321), .O(n469) );
  NR2T U858 ( .I1(n1112), .I2(n563), .O(n1095) );
  NR2T U859 ( .I1(n918), .I2(n513), .O(n908) );
  ND3 U860 ( .I1(n1061), .I2(n1062), .I3(n1063), .O(n1060) );
  AOI13HS U861 ( .B1(n539), .B2(n1078), .B3(n1079), .A1(n1080), .O(n1062) );
  OA22 U862 ( .A1(n1084), .A2(n46), .B1(n2397), .B2(n535), .O(n1061) );
  AOI112P U863 ( .C1(n46), .C2(n42), .A1(n1064), .B1(n1065), .O(n1063) );
  OAI112 U864 ( .C1(n1233), .C2(n2318), .A1(n1234), .B1(n1235), .O(n465) );
  ND2 U865 ( .I1(n1236), .I2(n1237), .O(n1234) );
  AOI13S U866 ( .B1(n485), .B2(n474), .B3(n1238), .A1(n1239), .O(n1233) );
  AOI112P U867 ( .C1(n1240), .C2(n1241), .A1(n485), .B1(n474), .O(n1239) );
  AOI112P U868 ( .C1(n2424), .C2(n112), .A1(n113), .B1(n114), .O(n110) );
  OAI112S U869 ( .C1(n135), .C2(n124), .A1(n136), .B1(n137), .O(n112) );
  MOAI1 U870 ( .A1(n115), .A2(n116), .B1(n2423), .B2(n118), .O(n114) );
  OAI112S U871 ( .C1(n2430), .C2(n131), .A1(n132), .B1(n133), .O(n113) );
  NR2T U872 ( .I1(n1054), .I2(n1042), .O(n1044) );
  NR2T U873 ( .I1(n539), .I2(n1083), .O(n1066) );
  ND3P U874 ( .I1(n388), .I2(n1817), .I3(n374), .O(n2270) );
  AOI13HS U875 ( .B1(n1749), .B2(n2377), .B3(n722), .A1(n1750), .O(n1748) );
  OAI12S U876 ( .B1(n2369), .B2(n725), .A1(n724), .O(n1749) );
  OA12 U877 ( .B1(n72), .B2(n1751), .A1(n2367), .O(n1750) );
  AOI12S U878 ( .B1(n2369), .B2(n715), .A1(n2377), .O(n1751) );
  NR2T U879 ( .I1(n2350), .I2(n582), .O(n591) );
  INV2 U880 ( .I(n1859), .O(n1029) );
  AOI13HS U881 ( .B1(n405), .B2(n131), .B3(n406), .A1(n135), .O(n404) );
  AOI13HS U882 ( .B1(n2427), .B2(n407), .B3(n138), .A1(n408), .O(n406) );
  NR2 U883 ( .I1(n409), .I2(n124), .O(n408) );
  NR2P U884 ( .I1(n46), .I2(n45), .O(n1076) );
  NR2T U885 ( .I1(n2354), .I2(n2356), .O(n695) );
  ND3P U886 ( .I1(n307), .I2(n850), .I3(n2338), .O(n1291) );
  NR2P U887 ( .I1(n518), .I2(n500), .O(n1261) );
  NR3P U888 ( .I1(n1850), .I2(n1851), .I3(n1852), .O(n1849) );
  OAI22 U889 ( .A1(n187), .A2(n1023), .B1(n585), .B2(n582), .O(n1852) );
  AO222 U890 ( .A1(n2351), .A2(n1854), .B1(n1030), .B2(n589), .C1(n582), .C2(
        n1855), .O(n1851) );
  OAI112S U891 ( .C1(n2351), .C2(n177), .A1(n584), .B1(n1011), .O(n1850) );
  ND2P U892 ( .I1(n338), .I2(n2331), .O(n335) );
  NR3P U893 ( .I1(n1903), .I2(n1904), .I3(n1905), .O(n1902) );
  OAI22 U894 ( .A1(n605), .A2(n608), .B1(n1049), .B2(n215), .O(n1905) );
  AO222 U895 ( .A1(n2346), .A2(n1907), .B1(n1055), .B2(n612), .C1(n605), .C2(
        n1908), .O(n1904) );
  OAI112S U896 ( .C1(n2346), .C2(n205), .A1(n607), .B1(n1036), .O(n1903) );
  ND3P U897 ( .I1(n146), .I2(n2415), .I3(n2414), .O(n1413) );
  NR3P U898 ( .I1(n663), .I2(n664), .I3(n665), .O(n662) );
  ND3 U899 ( .I1(n676), .I2(n677), .I3(n678), .O(n664) );
  MOAI1 U900 ( .A1(n666), .A2(n2353), .B1(n2353), .B2(n667), .O(n665) );
  OR3B2 U901 ( .I1(n106), .B1(n683), .B2(n684), .O(n663) );
  AO222 U902 ( .A1(n789), .A2(n1409), .B1(n1410), .B2(n1411), .C1(n788), .C2(
        n1412), .O(n461) );
  NR2 U903 ( .I1(n2409), .I2(n2406), .O(n1411) );
  NR2 U904 ( .I1(n1413), .I2(n2404), .O(n1410) );
  OAI12S U905 ( .B1(n2411), .B2(n790), .A1(n1414), .O(n1409) );
  NR3P U906 ( .I1(n765), .I2(n766), .I3(n767), .O(n764) );
  MOAI1 U907 ( .A1(n2411), .A2(n157), .B1(n457), .B2(n158), .O(n767) );
  OAI112S U908 ( .C1(n770), .C2(n2417), .A1(n771), .B1(n772), .O(n766) );
  OAI112S U909 ( .C1(n2408), .C2(n151), .A1(n780), .B1(n781), .O(n765) );
  NR3P U910 ( .I1(n733), .I2(n734), .I3(n735), .O(n732) );
  MOAI1 U911 ( .A1(n2428), .A2(n128), .B1(n426), .B2(n130), .O(n735) );
  OAI112S U912 ( .C1(n738), .C2(n2432), .A1(n739), .B1(n740), .O(n734) );
  OAI112S U913 ( .C1(n2423), .C2(n121), .A1(n748), .B1(n749), .O(n733) );
  BUF2 U914 ( .I(n150), .O(n2414) );
  NR2P U915 ( .I1(n332), .I2(n897), .O(n1332) );
  ND2P U916 ( .I1(n338), .I2(n334), .O(n330) );
  INV2 U917 ( .I(n2323), .O(n918) );
  AOI13HS U918 ( .B1(n357), .B2(n2218), .B3(n636), .A1(n2219), .O(n2211) );
  INV2 U919 ( .I(n638), .O(n2218) );
  NR3P U920 ( .I1(n637), .I2(n2315), .I3(n357), .O(n2219) );
  BUF2 U921 ( .I(n863), .O(n2340) );
  NR3P U922 ( .I1(n742), .I2(n1354), .I3(n135), .O(n1353) );
  ND3P U923 ( .I1(n186), .I2(n2351), .I3(n1853), .O(n1019) );
  AOI112P U924 ( .C1(n718), .C2(n65), .A1(n719), .B1(n720), .O(n717) );
  NR2 U925 ( .I1(n2375), .I2(n68), .O(n720) );
  ND3P U926 ( .I1(n282), .I2(n2388), .I3(n270), .O(n268) );
  NR2P U927 ( .I1(n862), .I2(n309), .O(n314) );
  OAI112 U928 ( .C1(n752), .C2(n753), .A1(n754), .B1(n755), .O(n429) );
  INV2 U929 ( .I(n758), .O(n753) );
  ND3 U930 ( .I1(n417), .I2(n129), .I3(n756), .O(n755) );
  ND3 U931 ( .I1(n2431), .I2(n2420), .I3(n757), .O(n754) );
  NR2T U932 ( .I1(n2356), .I2(n689), .O(n988) );
  ND3P U933 ( .I1(n2338), .I2(n867), .I3(n2343), .O(n1976) );
  OAI112 U934 ( .C1(n2069), .C2(n2070), .A1(n2071), .B1(n2072), .O(n1256) );
  INV2 U935 ( .I(n2066), .O(n2069) );
  ND3 U936 ( .I1(n1262), .I2(n500), .I3(n908), .O(n2071) );
  AOI13HS U937 ( .B1(n1261), .B2(n2330), .B3(n914), .A1(n2073), .O(n2072) );
  NR2T U938 ( .I1(n2368), .I2(n722), .O(n956) );
  OAI112 U939 ( .C1(n370), .C2(n2190), .A1(n2191), .B1(n2192), .O(n1183) );
  AO12 U940 ( .B1(n1190), .B2(n2195), .A1(n2196), .O(n2191) );
  OR3B2 U941 ( .I1(n2193), .B1(n352), .B2(n2194), .O(n2192) );
  ND2P U942 ( .I1(n1249), .I2(n485), .O(n488) );
  ND3P U943 ( .I1(n252), .I2(n254), .I3(n243), .O(n240) );
  OAI112 U944 ( .C1(n1563), .C2(n1559), .A1(n1564), .B1(n1565), .O(n1068) );
  ND3 U945 ( .I1(n1073), .I2(n2395), .I3(n43), .O(n1565) );
  ND3 U946 ( .I1(n1076), .I2(n44), .I3(n32), .O(n1564) );
  OA12 U947 ( .B1(n533), .B2(n36), .A1(n535), .O(n1563) );
  OAI112 U948 ( .C1(n1598), .C2(n1132), .A1(n1599), .B1(n1600), .O(n1128) );
  ND3 U949 ( .I1(n1602), .I2(n2393), .I3(n1603), .O(n1599) );
  AOI13HS U950 ( .B1(n1134), .B2(n254), .B3(n818), .A1(n1601), .O(n1600) );
  NR3P U951 ( .I1(n238), .I2(n815), .I3(n806), .O(n1601) );
  BUF2 U952 ( .I(n90), .O(n2363) );
  OAI112 U953 ( .C1(n1667), .C2(n1159), .A1(n1668), .B1(n1669), .O(n1155) );
  ND3 U954 ( .I1(n1673), .I2(n2382), .I3(n1674), .O(n1668) );
  AOI13HS U955 ( .B1(n1162), .B2(n270), .B3(n1670), .A1(n1671), .O(n1669) );
  NR3P U956 ( .I1(n1672), .I2(n840), .I3(n274), .O(n1671) );
  BUF2 U957 ( .I(n863), .O(n2339) );
  OAI12 U958 ( .B1(n2344), .B2(n1294), .A1(n308), .O(n313) );
  INV2 U959 ( .I(n1961), .O(n388) );
  ND3P U960 ( .I1(n2382), .I2(n282), .I3(n831), .O(n838) );
  BUF2 U961 ( .I(n150), .O(n2413) );
  NR2P U962 ( .I1(n862), .I2(n870), .O(n1301) );
  INV2 U963 ( .I(n2394), .O(n525) );
  NR2P U964 ( .I1(n2355), .I2(n990), .O(n672) );
  OA12 U965 ( .B1(n1485), .B2(n2402), .A1(n1486), .O(n546) );
  ND3 U966 ( .I1(n1105), .I2(n1487), .I3(n2402), .O(n1486) );
  OA12 U967 ( .B1(n1488), .B2(n558), .A1(n1489), .O(n1485) );
  MOAI1 U968 ( .A1(n558), .A2(n2400), .B1(n1110), .B2(n2400), .O(n1487) );
  OA12 U969 ( .B1(n1551), .B2(n2397), .A1(n1552), .O(n523) );
  OA12 U970 ( .B1(n1554), .B2(n534), .A1(n1555), .O(n1551) );
  ND3 U971 ( .I1(n1076), .I2(n1553), .I3(n2397), .O(n1552) );
  MOAI1 U972 ( .A1(n534), .A2(n2394), .B1(n1081), .B2(n2395), .O(n1553) );
  OAI112 U973 ( .C1(n228), .C2(n1914), .A1(n1915), .B1(n1916), .O(n596) );
  ND3 U974 ( .I1(n610), .I2(n1044), .I3(n1919), .O(n1915) );
  OA22 U975 ( .A1(n1917), .A2(n1040), .B1(n1043), .B2(n1045), .O(n1916) );
  OAI12 U976 ( .B1(n101), .B2(n2356), .A1(n690), .O(n670) );
  NR2P U977 ( .I1(n634), .I2(n627), .O(n1185) );
  OAI12 U978 ( .B1(n541), .B2(n37), .A1(n1077), .O(n42) );
  ND3 U979 ( .I1(n41), .I2(n44), .I3(n1071), .O(n1077) );
  BUF2 U980 ( .I(n74), .O(n2378) );
  BUF2 U981 ( .I(n348), .O(n2314) );
  OA222 U982 ( .A1(n2285), .A2(n2275), .B1(n2282), .B2(n2286), .C1(n2287), 
        .C2(n2270), .O(n643) );
  INV2 U983 ( .I(n1211), .O(n2287) );
  OA22 U984 ( .A1(n389), .A2(n2005), .B1(n388), .B2(n658), .O(n2286) );
  INV2 U985 ( .I(n1100), .O(n557) );
  ND2P U986 ( .I1(n1081), .I2(n525), .O(n536) );
  BUF2 U987 ( .I(n348), .O(n2315) );
  NR2P U988 ( .I1(n538), .I2(n1078), .O(n532) );
  OAI12 U989 ( .B1(n368), .B2(n634), .A1(n2217), .O(n628) );
  ND3 U990 ( .I1(n357), .I2(n634), .I3(n368), .O(n2217) );
  ND3 U991 ( .I1(n605), .I2(n603), .I3(n222), .O(n1914) );
  ND2P U992 ( .I1(n513), .I2(n2323), .O(n517) );
  BUF2 U993 ( .I(n90), .O(n2364) );
  NR2P U994 ( .I1(n562), .I2(n1107), .O(n556) );
  OAI112S U995 ( .C1(n468), .C2(n488), .A1(n475), .B1(n1242), .O(n2162) );
  OAI12 U996 ( .B1(n691), .B2(n692), .A1(n693), .O(n93) );
  INV2 U997 ( .I(n695), .O(n692) );
  OAI112S U998 ( .C1(n694), .C2(n672), .A1(n2353), .B1(n101), .O(n693) );
  NR2 U999 ( .I1(n2357), .I2(n674), .O(n694) );
  ND3 U1000 ( .I1(n198), .I2(n587), .I3(n1874), .O(n1868) );
  ND3 U1001 ( .I1(n2352), .I2(n1875), .I3(n591), .O(n1867) );
  AOI13HS U1002 ( .B1(n1024), .B2(n2351), .B3(n1865), .A1(n576), .O(n1869) );
  ND3 U1003 ( .I1(n357), .I2(n2315), .I3(n2194), .O(n2216) );
  INV2 U1004 ( .I(n1071), .O(n533) );
  ND3 U1005 ( .I1(n46), .I2(n44), .I3(n1078), .O(n1558) );
  ND2P U1006 ( .I1(n215), .I2(n603), .O(n1043) );
  ND3 U1007 ( .I1(n357), .I2(n2315), .I3(n359), .O(n2209) );
  ND3 U1008 ( .I1(n226), .I2(n610), .I3(n1927), .O(n1921) );
  ND3 U1009 ( .I1(n1928), .I2(n2349), .I3(n614), .O(n1920) );
  AOI13 U1010 ( .B1(n1050), .B2(n2346), .B3(n1918), .A1(n599), .O(n1922) );
  ND3 U1011 ( .I1(n512), .I2(n2083), .I3(n908), .O(n910) );
  BUF2 U1012 ( .I(n2171), .O(n2438) );
  BUF2 U1013 ( .I(n192), .O(n2352) );
  BUF2 U1014 ( .I(n92), .O(n2359) );
  INV2 U1015 ( .I(n1004), .O(n102) );
  INV2 U1016 ( .I(n972), .O(n75) );
  BUF2 U1017 ( .I(n117), .O(n2422) );
  MOAI1P U1018 ( .A1(n323), .A2(n2017), .B1(n1332), .B2(n2018), .O(n879) );
  OA22 U1019 ( .A1(n1318), .A2(n2019), .B1(n1316), .B2(n2021), .O(n2017) );
  OAI12S U1020 ( .B1(n2336), .B2(n2019), .A1(n2020), .O(n2018) );
  ND2P U1021 ( .I1(n605), .I2(n2347), .O(n227) );
  BUF2 U1022 ( .I(n2171), .O(n2439) );
  INV2 U1023 ( .I(n309), .O(n870) );
  ND3 U1024 ( .I1(n252), .I2(n806), .I3(n2392), .O(n1608) );
  OR3B2 U1025 ( .I1(n759), .B1(n116), .B2(n129), .O(n1359) );
  ND3 U1026 ( .I1(n2433), .I2(n419), .I3(n1363), .O(n1360) );
  BUF2 U1027 ( .I(n2172), .O(n2435) );
  BUF2 U1028 ( .I(n453), .O(n2411) );
  BUF2 U1029 ( .I(n421), .O(n2428) );
  NR2P U1030 ( .I1(n2422), .I2(n122), .O(n1367) );
  AO12 U1031 ( .B1(n400), .B2(n948), .A1(n401), .O(n61) );
  OAI22 U1032 ( .A1(n961), .A2(n75), .B1(n958), .B2(n702), .O(n400) );
  AN3 U1033 ( .I1(n957), .I2(n2376), .I3(n953), .O(n401) );
  MOAI1P U1034 ( .A1(n1870), .A2(n592), .B1(n1871), .B2(n1872), .O(n576) );
  OAI12S U1035 ( .B1(n187), .B2(n200), .A1(n1873), .O(n1872) );
  OA13 U1036 ( .B1(n1017), .B2(n176), .B3(n186), .A1(n1861), .O(n1870) );
  ND3 U1037 ( .I1(n187), .I2(n590), .I3(n1029), .O(n1873) );
  OAI12 U1038 ( .B1(n2379), .B2(n2368), .A1(n724), .O(n704) );
  OAI112S U1039 ( .C1(n2367), .C2(n963), .A1(n1752), .B1(n1753), .O(n1730) );
  MOAI1 U1040 ( .A1(n77), .A2(n1748), .B1(n966), .B2(n2371), .O(n1731) );
  ND3 U1041 ( .I1(n1754), .I2(n709), .I3(n718), .O(n1753) );
  OAI112S U1042 ( .C1(n2354), .C2(n995), .A1(n1814), .B1(n1815), .O(n1792) );
  MOAI1 U1043 ( .A1(n1810), .A2(n2361), .B1(n998), .B2(n2358), .O(n1793) );
  ND3 U1044 ( .I1(n1816), .I2(n674), .I3(n685), .O(n1815) );
  ND3 U1045 ( .I1(n819), .I2(n806), .I3(n1135), .O(n1129) );
  ND3 U1046 ( .I1(n817), .I2(n1134), .I3(n818), .O(n1130) );
  OA22 U1047 ( .A1(n811), .A2(n1132), .B1(n238), .B2(n1133), .O(n1131) );
  NR2P U1048 ( .I1(n680), .I2(n2355), .O(n1806) );
  NR2P U1049 ( .I1(n713), .I2(n2368), .O(n1744) );
  BUF2 U1050 ( .I(n369), .O(n2181) );
  OAI12S U1051 ( .B1(n2357), .B2(n101), .A1(n102), .O(n96) );
  MAOI1 U1052 ( .A1(n1330), .A2(n2026), .B1(n2027), .B2(n2028), .O(n321) );
  OAI12 U1053 ( .B1(n334), .B2(n335), .A1(n2024), .O(n2026) );
  OAI12S U1054 ( .B1(n2029), .B2(n2030), .A1(n323), .O(n2028) );
  INV2 U1055 ( .I(n1317), .O(n2030) );
  AO222 U1056 ( .A1(n1207), .A2(n1208), .B1(n1209), .B2(n1210), .C1(n1211), 
        .C2(n1212), .O(n642) );
  AO12 U1057 ( .B1(n380), .B2(n1213), .A1(n1214), .O(n1210) );
  OA12 U1058 ( .B1(n158), .B2(n1417), .A1(n1418), .O(n780) );
  ND3 U1059 ( .I1(n1419), .I2(n2416), .I3(n1420), .O(n1418) );
  AOI13HS U1060 ( .B1(n443), .B2(n439), .B3(n2414), .A1(n1421), .O(n1417) );
  NR2 U1061 ( .I1(n776), .I2(n2406), .O(n1420) );
  OAI12 U1062 ( .B1(n1003), .B2(n2363), .A1(n669), .O(n103) );
  AOI12S U1063 ( .B1(n672), .B2(n101), .A1(n1005), .O(n1003) );
  NR2P U1064 ( .I1(n517), .I2(n500), .O(n2062) );
  OA112 U1065 ( .C1(n2144), .C2(n485), .A1(n2145), .B1(n2146), .O(n1235) );
  ND3 U1066 ( .I1(n2147), .I2(n2319), .I3(n1238), .O(n2146) );
  ND3 U1067 ( .I1(n2317), .I2(n2148), .I3(n1237), .O(n2145) );
  OA112 U1068 ( .C1(n1598), .C2(n1133), .A1(n1126), .B1(n1604), .O(n249) );
  OA222 U1069 ( .A1(n238), .A2(n1132), .B1(n1605), .B2(n1606), .C1(n240), .C2(
        n1607), .O(n1604) );
  ND3 U1070 ( .I1(n236), .I2(n806), .I3(n809), .O(n1605) );
  ND2 U1071 ( .I1(n817), .I2(n1602), .O(n1606) );
  OA112 U1072 ( .C1(n1667), .C2(n1160), .A1(n1153), .B1(n1675), .O(n277) );
  OA222 U1073 ( .A1(n266), .A2(n1159), .B1(n1676), .B2(n1677), .C1(n268), .C2(
        n1678), .O(n1675) );
  ND2 U1074 ( .I1(n1161), .I2(n2380), .O(n1678) );
  ND3 U1075 ( .I1(n2390), .I2(n2384), .I3(n831), .O(n1676) );
  OA112 U1076 ( .C1(n834), .C2(n1160), .A1(n1683), .B1(n1684), .O(n1154) );
  ND3 U1077 ( .I1(n270), .I2(n842), .I3(n1162), .O(n1683) );
  AOI13HS U1078 ( .B1(n840), .B2(n1670), .B3(n841), .A1(n1685), .O(n1684) );
  NR3P U1079 ( .I1(n1679), .I2(n840), .I3(n274), .O(n1685) );
  INV2 U1080 ( .I(n341), .O(n1316) );
  INV2 U1081 ( .I(n2194), .O(n637) );
  OAI112S U1082 ( .C1(n2165), .C2(n2164), .A1(n2166), .B1(n927), .O(n2160) );
  INV2 U1083 ( .I(n1249), .O(n2165) );
  ND3 U1084 ( .I1(n2164), .I2(n2318), .I3(n2167), .O(n2166) );
  NR2 U1085 ( .I1(n484), .I2(n485), .O(n2167) );
  AO222 U1086 ( .A1(n485), .A2(n2140), .B1(n2141), .B2(n2142), .C1(n2143), 
        .C2(n1237), .O(n1232) );
  NR2 U1087 ( .I1(n2317), .I2(n485), .O(n2141) );
  AO22 U1088 ( .A1(n932), .A2(n1236), .B1(n2143), .B2(n934), .O(n2140) );
  ND2P U1089 ( .I1(encrypt_shift[1]), .I2(encrypt_shift[0]), .O(n2090) );
  AO222 U1090 ( .A1(n2059), .A2(n2326), .B1(n2060), .B2(n2061), .C1(n2062), 
        .C2(n1262), .O(n1257) );
  NR2 U1091 ( .I1(n513), .I2(n2328), .O(n2060) );
  AO22 U1092 ( .A1(n912), .A2(n1261), .B1(n2062), .B2(n914), .O(n2059) );
  INV2 U1093 ( .I(n1221), .O(n645) );
  OAI12S U1094 ( .B1(n1964), .B2(n309), .A1(n1965), .O(n1962) );
  AOI13HS U1095 ( .B1(n2340), .B2(n1294), .B3(n305), .A1(n1968), .O(n1964) );
  ND3 U1096 ( .I1(n309), .I2(n869), .I3(n2341), .O(n1965) );
  NR2 U1097 ( .I1(n1969), .I2(n850), .O(n1968) );
  INV2 U1098 ( .I(n774), .O(n153) );
  ND3 U1099 ( .I1(n2276), .I2(n380), .I3(n1221), .O(n2284) );
  AO222 U1100 ( .A1(n1074), .A2(n1556), .B1(n1557), .B2(n1078), .C1(n1067), 
        .C2(n1081), .O(n1065) );
  NR2 U1101 ( .I1(n534), .I2(n1559), .O(n1557) );
  OAI12S U1102 ( .B1(n2396), .B2(n533), .A1(n37), .O(n1556) );
  ND3 U1103 ( .I1(n982), .I2(n983), .I3(n984), .O(n686) );
  ND3 U1104 ( .I1(n992), .I2(n2360), .I3(n695), .O(n982) );
  AOI13HS U1105 ( .B1(n101), .B2(n985), .B3(n986), .A1(n987), .O(n984) );
  ND3 U1106 ( .I1(n2354), .I2(n2356), .I3(n991), .O(n983) );
  NR2P U1107 ( .I1(n541), .I2(n533), .O(n1543) );
  ND3 U1108 ( .I1(n2384), .I2(n2387), .I3(n2382), .O(n1679) );
  INV2 U1109 ( .I(n2200), .O(n370) );
  ND3 U1110 ( .I1(n352), .I2(n2200), .I3(n1197), .O(n2208) );
  OAI12S U1111 ( .B1(n62), .B2(n63), .A1(n64), .O(n60) );
  ND3 U1112 ( .I1(n65), .I2(n2374), .I3(n62), .O(n64) );
  OA12 U1113 ( .B1(n2366), .B2(n67), .A1(n68), .O(n63) );
  MAOI1 U1114 ( .A1(n69), .A2(n2372), .B1(n70), .B2(n2373), .O(n67) );
  OAI12S U1115 ( .B1(n468), .B2(n488), .A1(n936), .O(n933) );
  NR2 U1116 ( .I1(n938), .I2(n2321), .O(n931) );
  INV2 U1117 ( .I(n469), .O(n935) );
  OAI12S U1118 ( .B1(n2324), .B2(n516), .A1(n917), .O(n913) );
  NR2 U1119 ( .I1(n2330), .I2(n919), .O(n911) );
  INV2 U1120 ( .I(n497), .O(n915) );
  NR2P U1121 ( .I1(n645), .I2(n1961), .O(n2271) );
  ND2P U1122 ( .I1(encrypt_shift[1]), .I2(n2311), .O(n2092) );
  NR2P U1123 ( .I1(n565), .I2(n557), .O(n1477) );
  AO222 U1124 ( .A1(n2315), .A2(n2201), .B1(n2202), .B2(n2203), .C1(n1189), 
        .C2(n2204), .O(n1182) );
  NR2 U1125 ( .I1(n359), .I2(n357), .O(n2203) );
  INV2 U1126 ( .I(n1190), .O(n2204) );
  OAI12S U1127 ( .B1(n2206), .B2(n2207), .A1(n2208), .O(n2201) );
  ND2P U1128 ( .I1(encrypt_shift[0]), .I2(n2312), .O(n2094) );
  AO222 U1129 ( .A1(n2277), .A2(n2005), .B1(n2278), .B2(n2279), .C1(n1212), 
        .C2(n1214), .O(n1205) );
  NR2 U1130 ( .I1(n1802), .I2(n1961), .O(n2278) );
  OAI12S U1131 ( .B1(n2282), .B2(n2283), .A1(n2284), .O(n2277) );
  NR2 U1132 ( .I1(n374), .I2(n2275), .O(n2279) );
  ND3 U1133 ( .I1(n950), .I2(n951), .I3(n952), .O(n719) );
  ND3 U1134 ( .I1(n960), .I2(n2373), .I3(n729), .O(n950) );
  AOI13HS U1135 ( .B1(n2379), .B2(n953), .B3(n954), .A1(n955), .O(n952) );
  ND3 U1136 ( .I1(n2369), .I2(n2367), .I3(n959), .O(n951) );
  ND3 U1137 ( .I1(n43), .I2(n2395), .I3(n1081), .O(n1555) );
  ND2P U1138 ( .I1(n1332), .I2(n2334), .O(n2025) );
  ND3 U1139 ( .I1(n729), .I2(n2376), .I3(n1736), .O(n1734) );
  NR2P U1140 ( .I1(n2021), .I2(n2336), .O(n1315) );
  AO222 U1141 ( .A1(n2340), .A2(n1286), .B1(n1287), .B2(n1288), .C1(n855), 
        .C2(n1289), .O(n853) );
  NR2 U1143 ( .I1(n1290), .I2(n2339), .O(n1287) );
  OAI12S U1144 ( .B1(n1291), .B2(n1292), .A1(n1293), .O(n1286) );
  OR3 U1145 ( .I1(n303), .I2(n1294), .I3(n1290), .O(n1293) );
  AO222 U1146 ( .A1(n1313), .A2(n2334), .B1(n1314), .B2(n323), .C1(n882), .C2(
        n1315), .O(n880) );
  NR2 U1147 ( .I1(n1316), .I2(n1317), .O(n1314) );
  OAI12S U1148 ( .B1(n1317), .B2(n1318), .A1(n1319), .O(n1313) );
  OR3 U1149 ( .I1(n330), .I2(n1316), .I3(n2332), .O(n1319) );
  INV2 U1150 ( .I(n122), .O(n125) );
  INV2 U1151 ( .I(n224), .O(n228) );
  ND3 U1152 ( .I1(n2414), .I2(n2405), .I3(n788), .O(n785) );
  MOAI1 U1153 ( .A1(n1864), .A2(n1029), .B1(n580), .B2(n1018), .O(n1875) );
  INV2 U1154 ( .I(n1213), .O(n658) );
  AO222 U1155 ( .A1(n323), .A2(n2031), .B1(n2032), .B2(n1330), .C1(n2033), 
        .C2(n2029), .O(n884) );
  INV2 U1156 ( .I(n2025), .O(n2033) );
  NR2 U1157 ( .I1(n2331), .I2(n329), .O(n2032) );
  MOAI1 U1158 ( .A1(n2019), .A2(n1316), .B1(n1327), .B2(n2029), .O(n2031) );
  OA12 U1159 ( .B1(n1980), .B2(n1981), .A1(n1982), .O(n294) );
  AOI12S U1160 ( .B1(n1307), .B2(n867), .A1(n856), .O(n1980) );
  OAI112S U1161 ( .C1(n1983), .C2(n1288), .A1(n2341), .B1(n855), .O(n1982) );
  ND2 U1162 ( .I1(n1918), .I2(n204), .O(n1040) );
  ND2 U1163 ( .I1(n538), .I2(n46), .O(n1554) );
  INV2 U1164 ( .I(n1670), .O(n266) );
  INV2 U1165 ( .I(n842), .O(n1667) );
  AO222 U1166 ( .A1(n62), .A2(n1745), .B1(n1746), .B2(n1747), .C1(n959), .C2(
        n956), .O(n949) );
  NR2 U1167 ( .I1(n722), .I2(n2371), .O(n1747) );
  NR2 U1168 ( .I1(n2372), .I2(n1737), .O(n1746) );
  AO22 U1169 ( .A1(n1744), .A2(n972), .B1(n1736), .B2(n729), .O(n1745) );
  INV2 U1170 ( .I(n668), .O(n673) );
  INV2 U1171 ( .I(n1379), .O(n2490) );
  INV2 U1172 ( .I(n41), .O(n36) );
  ND3 U1173 ( .I1(n975), .I2(n976), .I3(n977), .O(n974) );
  NR2 U1174 ( .I1(n997), .I2(n998), .O(n976) );
  AOI13HS U1175 ( .B1(n2360), .B2(n103), .B3(n689), .A1(n999), .O(n975) );
  AOI112P U1176 ( .C1(n2353), .C2(n978), .A1(n979), .B1(n107), .O(n977) );
  AO222 U1177 ( .A1(n2364), .A2(n1807), .B1(n1808), .B2(n1809), .C1(n991), 
        .C2(n988), .O(n981) );
  NR2 U1178 ( .I1(n2358), .I2(n689), .O(n1809) );
  NR2 U1179 ( .I1(n1799), .I2(n2359), .O(n1808) );
  AO22 U1180 ( .A1(n1806), .A2(n1004), .B1(n1798), .B2(n695), .O(n1807) );
  ND3 U1181 ( .I1(n922), .I2(n923), .I3(n924), .O(n921) );
  NR2 U1182 ( .I1(n939), .I2(n465), .O(n922) );
  OA222 U1183 ( .A1(n925), .A2(n471), .B1(n926), .B2(n485), .C1(n473), .C2(
        n927), .O(n924) );
  OA13 U1184 ( .B1(n473), .B2(n928), .B3(n929), .A1(n930), .O(n926) );
  OA12 U1185 ( .B1(n1609), .B2(n243), .A1(n1610), .O(n1126) );
  ND3 U1186 ( .I1(n809), .I2(n1611), .I3(n1147), .O(n1610) );
  OA22 U1187 ( .A1(n815), .A2(n811), .B1(n248), .B2(n238), .O(n1609) );
  MOAI1 U1188 ( .A1(n1598), .A2(n2393), .B1(n2393), .B2(n1134), .O(n1611) );
  OA222 U1189 ( .A1(n252), .A2(n253), .B1(n254), .B2(n255), .C1(n256), .C2(
        n257), .O(n251) );
  INV2 U1190 ( .I(n258), .O(n256) );
  OA12 U1191 ( .B1(n270), .B2(n1680), .A1(n1681), .O(n1153) );
  ND3 U1192 ( .I1(n831), .I2(n1682), .I3(n1174), .O(n1681) );
  OA22 U1193 ( .A1(n838), .A2(n834), .B1(n276), .B2(n266), .O(n1680) );
  MOAI1 U1194 ( .A1(n1667), .A2(n2381), .B1(n2381), .B2(n1161), .O(n1682) );
  ND3 U1195 ( .I1(n943), .I2(n944), .I3(n945), .O(n942) );
  NR2 U1196 ( .I1(n965), .I2(n966), .O(n944) );
  AOI13HS U1197 ( .B1(n76), .B2(n2373), .B3(n722), .A1(n967), .O(n943) );
  AOI112P U1198 ( .C1(n946), .C2(n2366), .A1(n947), .B1(n80), .O(n945) );
  OA222 U1199 ( .A1(n2387), .A2(n281), .B1(n282), .B2(n283), .C1(n284), .C2(
        n285), .O(n279) );
  INV2 U1200 ( .I(n286), .O(n284) );
  NR2P U1201 ( .I1(n920), .I2(n1256), .O(n494) );
  ND3 U1202 ( .I1(n1090), .I2(n1091), .I3(n1092), .O(n1089) );
  AOI13HS U1203 ( .B1(n1107), .B2(n563), .B3(n1108), .A1(n1109), .O(n1091) );
  OA22 U1204 ( .A1(n551), .A2(n1113), .B1(n2401), .B2(n559), .O(n1090) );
  AOI112P U1205 ( .C1(n551), .C2(n19), .A1(n1093), .B1(n1094), .O(n1092) );
  ND3 U1206 ( .I1(n1595), .I2(n1596), .I3(n1597), .O(n1594) );
  MAOI1 U1207 ( .A1(n802), .A2(n814), .B1(n809), .B2(n816), .O(n1595) );
  AOI112P U1208 ( .C1(n806), .C2(n1619), .A1(n1620), .B1(n1141), .O(n1596) );
  AOI112P U1209 ( .C1(n258), .C2(n257), .A1(n803), .B1(n1128), .O(n1597) );
  INV2 U1210 ( .I(n912), .O(n506) );
  ND2 U1211 ( .I1(n1616), .I2(n1617), .O(n258) );
  ND3 U1212 ( .I1(n801), .I2(n2392), .I3(n1603), .O(n1617) );
  ND3 U1213 ( .I1(n1618), .I2(n814), .I3(n243), .O(n1616) );
  INV2 U1214 ( .I(n18), .O(n13) );
  AO222 U1215 ( .A1(n758), .A2(n1340), .B1(n1341), .B2(n1342), .C1(n757), .C2(
        n1343), .O(n430) );
  NR2 U1216 ( .I1(n2426), .I2(n2422), .O(n1342) );
  NR2 U1217 ( .I1(n1344), .I2(n2420), .O(n1341) );
  OAI12S U1218 ( .B1(n2428), .B2(n759), .A1(n1345), .O(n1340) );
  ND2 U1219 ( .I1(n562), .I2(n551), .O(n1488) );
  AN3 U1220 ( .I1(n1306), .I2(n867), .I3(n1307), .O(n315) );
  INV2 U1221 ( .I(n543), .O(n51) );
  INV2 U1223 ( .I(n567), .O(n27) );
  INV2 U1224 ( .I(n1327), .O(n1318) );
  OAI12S U1225 ( .B1(n89), .B2(n2363), .A1(n91), .O(n87) );
  ND3 U1226 ( .I1(n2360), .I2(n93), .I3(n2364), .O(n91) );
  OA12 U1227 ( .B1(n2353), .B2(n94), .A1(n95), .O(n89) );
  MAOI1 U1228 ( .A1(n2359), .A2(n96), .B1(n97), .B2(n2360), .O(n94) );
  OA112 U1229 ( .C1(n1318), .C2(n2020), .A1(n2022), .B1(n2023), .O(n878) );
  ND3 U1230 ( .I1(n1332), .I2(n323), .I3(n883), .O(n2023) );
  AO12 U1231 ( .B1(n1317), .B2(n2021), .A1(n2025), .O(n2022) );
  OA222 U1232 ( .A1(n361), .A2(n363), .B1(n364), .B2(n365), .C1(n366), .C2(
        n367), .O(n356) );
  ND2 U1233 ( .I1(n368), .I2(n366), .O(n365) );
  ND2 U1234 ( .I1(n2280), .I2(n370), .O(n364) );
  AN3 U1235 ( .I1(n1876), .I2(n1877), .I3(n1878), .O(n584) );
  ND3 U1236 ( .I1(n1016), .I2(n589), .I3(n591), .O(n1877) );
  OR3B2 U1237 ( .I1(n1019), .B1(n2352), .B2(n580), .O(n1876) );
  AOI13HS U1238 ( .B1(n1871), .B2(n1859), .B3(n1024), .A1(n1879), .O(n1878) );
  INV2 U1239 ( .I(n1208), .O(n2283) );
  OA22 U1240 ( .A1(n185), .A2(n186), .B1(n187), .B2(n188), .O(n184) );
  AOI13HS U1241 ( .B1(n187), .B2(n189), .B3(n176), .A1(n190), .O(n185) );
  NR2 U1242 ( .I1(n191), .I2(n192), .O(n190) );
  MAOI1 U1243 ( .A1(n193), .A2(n194), .B1(n195), .B2(n176), .O(n191) );
  OR2 U1244 ( .I1(n1608), .I2(n254), .O(n1132) );
  OR2 U1245 ( .I1(n1679), .I2(n282), .O(n1159) );
  OA22 U1246 ( .A1(n1139), .A2(n254), .B1(n806), .B2(n245), .O(n1138) );
  AOI12S U1247 ( .B1(n809), .B2(n1140), .A1(n1141), .O(n1139) );
  OAI12S U1248 ( .B1(n243), .B2(n1142), .A1(n239), .O(n1140) );
  AN3 U1249 ( .I1(n1426), .I2(n1427), .I3(n1428), .O(n782) );
  OR3B2 U1250 ( .I1(n790), .B1(n146), .B2(n159), .O(n1426) );
  ND3 U1251 ( .I1(n2418), .I2(n451), .I3(n1430), .O(n1427) );
  AOI13HS U1252 ( .B1(n158), .B2(n2414), .B3(n788), .A1(n1429), .O(n1428) );
  OA12 U1253 ( .B1(n743), .B2(n116), .A1(n137), .O(n738) );
  OA222 U1254 ( .A1(n2425), .A2(n744), .B1(n2421), .B2(n745), .C1(n135), .C2(
        n746), .O(n743) );
  ND2 U1255 ( .I1(n747), .I2(n122), .O(n745) );
  XNR2 U1256 ( .I1(n2425), .I2(n135), .O(n747) );
  OA222 U1257 ( .A1(n248), .A2(n257), .B1(n246), .B2(n815), .C1(n254), .C2(
        n239), .O(n805) );
  INV2 U1258 ( .I(n1344), .O(n1352) );
  INV2 U1259 ( .I(n882), .O(n2027) );
  ND3 U1260 ( .I1(n412), .I2(n413), .I3(n414), .O(n403) );
  ND3 U1261 ( .I1(n2427), .I2(n417), .I3(n418), .O(n413) );
  ND3 U1262 ( .I1(n2425), .I2(n415), .I3(n416), .O(n414) );
  OR3B2 U1263 ( .I1(n420), .B1(n2429), .B2(n422), .O(n412) );
  OA222 U1264 ( .A1(n22), .A2(n560), .B1(n561), .B2(n2402), .C1(n562), .C2(n14), .O(n550) );
  AOI112P U1265 ( .C1(n563), .C2(n18), .A1(n9), .B1(n564), .O(n561) );
  NR2 U1266 ( .I1(n17), .I2(n565), .O(n564) );
  INV2 U1267 ( .I(n1640), .O(n1375) );
  INV2 U1268 ( .I(encrypt_shift[0]), .O(n2311) );
  INV2 U1269 ( .I(n1642), .O(n1377) );
  INV2 U1270 ( .I(encrypt_shift[1]), .O(n2312) );
  ND2 U1271 ( .I1(n482), .I2(n483), .O(n477) );
  XNR2 U1272 ( .I1(n484), .I2(n474), .O(n482) );
  NR2 U1273 ( .I1(n594), .I2(n595), .O(n593) );
  ND3 U1274 ( .I1(n608), .I2(n205), .I3(n609), .O(n594) );
  OR3B2 U1275 ( .I1(n596), .B1(n206), .B2(n597), .O(n595) );
  AOI13HS U1276 ( .B1(n605), .B2(n217), .B3(n610), .A1(n611), .O(n609) );
  NR2 U1277 ( .I1(n619), .I2(n620), .O(n618) );
  OAI112S U1278 ( .C1(n623), .C2(n624), .A1(n625), .B1(n626), .O(n619) );
  OR3B2 U1279 ( .I1(n621), .B1(n351), .B2(n622), .O(n620) );
  OA22 U1280 ( .A1(n636), .A2(n637), .B1(n638), .B2(n635), .O(n623) );
  NR2 U1281 ( .I1(n640), .I2(n641), .O(n639) );
  OAI112S U1282 ( .C1(n644), .C2(n645), .A1(n646), .B1(n647), .O(n640) );
  OR3B2 U1283 ( .I1(n642), .B1(n395), .B2(n643), .O(n641) );
  OA22 U1284 ( .A1(n657), .A2(n658), .B1(n659), .B2(n656), .O(n644) );
  OAI112 U1285 ( .C1(n1497), .C2(n1493), .A1(n1498), .B1(n1499), .O(n1097) );
  ND3 U1286 ( .I1(n1102), .I2(n2400), .I3(n20), .O(n1499) );
  ND3 U1287 ( .I1(n1105), .I2(n21), .I3(n9), .O(n1498) );
  OA12 U1288 ( .B1(n557), .B2(n13), .A1(n559), .O(n1497) );
  NR2 U1289 ( .I1(n1180), .I2(n1181), .O(n1179) );
  ND3 U1290 ( .I1(n1191), .I2(n1192), .I3(n1193), .O(n1180) );
  OR3B2 U1291 ( .I1(n1182), .B1(n350), .B2(n622), .O(n1181) );
  OR3B2 U1292 ( .I1(n363), .B1(n1197), .B2(n634), .O(n1192) );
  ND3 U1293 ( .I1(n1560), .I2(n1561), .I3(n1562), .O(n542) );
  ND3 U1294 ( .I1(n1082), .I2(n1066), .I3(n538), .O(n1560) );
  ND3 U1295 ( .I1(n525), .I2(n1073), .I3(n1076), .O(n1561) );
  OA22 U1296 ( .A1(n44), .A2(n1555), .B1(n533), .B2(n1558), .O(n1562) );
  NR2 U1297 ( .I1(n317), .I2(n318), .O(n316) );
  OAI112S U1298 ( .C1(n323), .C2(n324), .A1(n325), .B1(n326), .O(n317) );
  OAI112S U1299 ( .C1(n319), .C2(n320), .A1(n321), .B1(n322), .O(n318) );
  ND3 U1300 ( .I1(n332), .I2(n333), .I3(n323), .O(n325) );
  NR2 U1301 ( .I1(n1124), .I2(n1125), .O(n1123) );
  OAI112S U1302 ( .C1(n1136), .C2(n801), .A1(n1137), .B1(n1138), .O(n1124) );
  ND3 U1303 ( .I1(n250), .I2(n1126), .I3(n1127), .O(n1125) );
  ND3 U1304 ( .I1(n252), .I2(n1143), .I3(n801), .O(n1137) );
  OA22 U1305 ( .A1(n1194), .A2(n359), .B1(n632), .B2(n367), .O(n1193) );
  AOI13HS U1306 ( .B1(n632), .B2(n635), .B3(n1185), .A1(n1195), .O(n1194) );
  NR3P U1307 ( .I1(n1196), .I2(n638), .I3(n368), .O(n1195) );
  XNR2 U1308 ( .I1(n357), .I2(n2181), .O(n1196) );
  NR2 U1309 ( .I1(n2138), .I2(n2139), .O(n2137) );
  AO222 U1310 ( .A1(n2316), .A2(n2160), .B1(n485), .B2(n2161), .C1(n474), .C2(
        n2162), .O(n2138) );
  ND3 U1311 ( .I1(n466), .I2(n1235), .I3(n923), .O(n2139) );
  OAI12S U1312 ( .B1(n471), .B2(n929), .A1(n930), .O(n2161) );
  NR2 U1313 ( .I1(n1406), .I2(n1407), .O(n1405) );
  OAI112S U1314 ( .C1(n1431), .C2(n2415), .A1(n1432), .B1(n1433), .O(n1406) );
  OAI112S U1315 ( .C1(n452), .C2(n442), .A1(n782), .B1(n1408), .O(n1407) );
  OA13 U1316 ( .B1(n455), .B2(n2410), .B3(n792), .A1(n437), .O(n1431) );
  NR2 U1317 ( .I1(n1009), .I2(n1010), .O(n1008) );
  AO2222 U1318 ( .A1(n580), .A2(n1020), .B1(n1021), .B2(n2351), .C1(n198), 
        .C2(n589), .D1(n187), .D2(n1022), .O(n1009) );
  OAI112S U1319 ( .C1(n2351), .C2(n183), .A1(n583), .B1(n1011), .O(n1010) );
  INV2 U1320 ( .I(n577), .O(n1021) );
  NR2 U1321 ( .I1(n202), .I2(n203), .O(n201) );
  OAI112S U1322 ( .C1(n209), .C2(n210), .A1(n211), .B1(n212), .O(n202) );
  OAI112S U1323 ( .C1(n204), .C2(n205), .A1(n206), .B1(n207), .O(n203) );
  INV2 U1324 ( .I(n222), .O(n210) );
  NR3P U1325 ( .I1(n879), .I2(n880), .I3(n881), .O(n322) );
  AO13 U1326 ( .B1(n882), .B2(n323), .B3(n883), .A1(n884), .O(n881) );
  ND2 U1327 ( .I1(n932), .I2(n471), .O(n1241) );
  NR2 U1328 ( .I1(n1229), .I2(n1230), .O(n1228) );
  OAI112S U1329 ( .C1(n474), .C2(n1242), .A1(n1243), .B1(n1244), .O(n1229) );
  OR3 U1330 ( .I1(n1231), .I2(n465), .I3(n1232), .O(n1230) );
  ND2 U1331 ( .I1(n473), .I2(n1250), .O(n1243) );
  NR2 U1332 ( .I1(n1309), .I2(n1310), .O(n1308) );
  OAI112S U1333 ( .C1(n1322), .C2(n2335), .A1(n1323), .B1(n1324), .O(n1309) );
  AO112 U1334 ( .C1(n332), .C2(n1311), .A1(n880), .B1(n1312), .O(n1310) );
  AOI13HS U1335 ( .B1(n892), .B2(n1325), .B3(n1326), .A1(n328), .O(n1324) );
  AN2 U1336 ( .I1(n606), .I2(n607), .O(n206) );
  AN3B1 U1337 ( .I1(n589), .I2(n590), .B1(n591), .O(n588) );
  AN3 U1338 ( .I1(n1865), .I2(n590), .I3(n587), .O(n1879) );
  INV2 U1339 ( .I(n485), .O(n480) );
  OR3B2 U1340 ( .I1(n465), .B1(n466), .B2(n467), .O(n464) );
  OA222 U1341 ( .A1(n468), .A2(n469), .B1(n470), .B2(n471), .C1(n472), .C2(
        n473), .O(n467) );
  OA222 U1342 ( .A1(n2317), .A2(n488), .B1(n489), .B2(n490), .C1(n478), .C2(
        n491), .O(n470) );
  OA222 U1343 ( .A1(n474), .A2(n475), .B1(n476), .B2(n477), .C1(n478), .C2(
        n479), .O(n472) );
  NR3P U1344 ( .I1(n697), .I2(n698), .I3(n699), .O(n696) );
  ND3 U1345 ( .I1(n710), .I2(n711), .I3(n712), .O(n698) );
  MOAI1 U1346 ( .A1(n700), .A2(n2366), .B1(n701), .B2(n2366), .O(n699) );
  OR3B2 U1347 ( .I1(n79), .B1(n716), .B2(n717), .O(n697) );
  INV2 U1348 ( .I(n44), .O(n529) );
  NR2 U1349 ( .I1(n2403), .I2(n1425), .O(n1424) );
  NR2 U1350 ( .I1(n575), .I2(n576), .O(n574) );
  AOI13HS U1351 ( .B1(n577), .B2(n188), .B3(n578), .A1(n2351), .O(n575) );
  ND3 U1352 ( .I1(n580), .I2(n193), .I3(n581), .O(n578) );
  NR2 U1353 ( .I1(n582), .I2(n2352), .O(n581) );
  OA112 U1354 ( .C1(n1012), .C2(n187), .A1(n1013), .B1(n1014), .O(n583) );
  OR3B2 U1355 ( .I1(n1017), .B1(n1018), .B2(n591), .O(n1013) );
  OA22 U1356 ( .A1(n590), .A2(n1015), .B1(n2352), .B2(n1019), .O(n1012) );
  OR3 U1357 ( .I1(n1015), .I2(n580), .I3(n1016), .O(n1014) );
  INV2 U1358 ( .I(n21), .O(n553) );
  INV2 U1359 ( .I(n135), .O(n120) );
  ND2 U1360 ( .I1(n546), .I2(n567), .O(n1093) );
  ND2 U1361 ( .I1(n523), .I2(n543), .O(n1064) );
  INV1 U1362 ( .I(n474), .O(n487) );
  INV2 U1363 ( .I(n850), .O(n311) );
  AN3 U1364 ( .I1(n2143), .I2(n485), .I3(n932), .O(n2154) );
  OR2 U1365 ( .I1(n432), .I2(n433), .O(n1959) );
  AO112 U1366 ( .C1(n850), .C2(n1971), .A1(n1285), .B1(n852), .O(n432) );
  AO112 U1367 ( .C1(n307), .C2(n1962), .A1(n1963), .B1(n871), .O(n433) );
  AO12 U1368 ( .B1(n103), .B2(n2362), .A1(n105), .O(n86) );
  AO12 U1369 ( .B1(n76), .B2(n77), .A1(n78), .O(n58) );
  AN3 U1370 ( .I1(n2062), .I2(n2327), .I3(n912), .O(n2073) );
  OA12 U1371 ( .B1(n254), .B2(n810), .A1(n253), .O(n808) );
  OA12 U1372 ( .B1(n243), .B2(n811), .A1(n812), .O(n810) );
  ND3 U1373 ( .I1(n801), .I2(n2393), .I3(n243), .O(n812) );
  ND2 U1374 ( .I1(n510), .I2(n511), .O(n505) );
  XNR2 U1375 ( .I1(n512), .I2(n513), .O(n510) );
  AOI112P U1376 ( .C1(n959), .C2(n948), .A1(n61), .B1(n1732), .O(n716) );
  AO13 U1377 ( .B1(n77), .B2(n956), .B3(n960), .A1(n1733), .O(n1732) );
  ND2 U1378 ( .I1(n1734), .I2(n1735), .O(n1733) );
  ND3 U1379 ( .I1(n62), .I2(n953), .I3(n972), .O(n1735) );
  OAI12 U1380 ( .B1(n1966), .B2(n305), .A1(n1967), .O(n869) );
  ND3 U1381 ( .I1(n850), .I2(n1294), .I3(n305), .O(n1967) );
  INV2 U1382 ( .I(n313), .O(n1966) );
  MOAI1 U1383 ( .A1(n257), .A2(n236), .B1(n806), .B2(n1142), .O(n1148) );
  INV2 U1384 ( .I(n244), .O(n1149) );
  OR2 U1385 ( .I1(n1373), .I2(n1440), .O(n399) );
  AO112 U1386 ( .C1(n426), .C2(n2421), .A1(n428), .B1(n429), .O(n1373) );
  AO112 U1387 ( .C1(n402), .C2(n2423), .A1(n403), .B1(n404), .O(n1440) );
  ND2 U1388 ( .I1(n1134), .I2(n2391), .O(n1607) );
  INV2 U1389 ( .I(n2356), .O(n100) );
  INV2 U1390 ( .I(n2369), .O(n73) );
  INV2 U1391 ( .I(n2416), .O(n164) );
  INV2 U1392 ( .I(n2382), .O(n264) );
  OR2 U1393 ( .I1(n14), .I2(n2400), .O(n1118) );
  XNR2 U1394 ( .I1(n1054), .I2(n2349), .O(n225) );
  NR3P U1395 ( .I1(n2395), .I2(n1083), .I3(n1087), .O(n47) );
  XNR2 U1396 ( .I1(n2412), .I2(n2404), .O(n163) );
  XNR2 U1397 ( .I1(n862), .I2(n867), .O(n865) );
  XNR2 U1398 ( .I1(n334), .I2(n2332), .O(n1329) );
  ND3P U1399 ( .I1(n146), .I2(n2405), .I3(n2418), .O(n442) );
  XNR2 U1400 ( .I1(n867), .I2(n2338), .O(n1303) );
  XNR2 U1401 ( .I1(n334), .I2(n332), .O(n892) );
  ND3P U1402 ( .I1(n275), .I2(n2381), .I3(n1174), .O(n281) );
  ND3P U1403 ( .I1(n247), .I2(n2393), .I3(n1147), .O(n253) );
  ND3P U1404 ( .I1(n101), .I2(n988), .I3(n1803), .O(n677) );
  ND3P U1405 ( .I1(n605), .I2(n1042), .I3(n612), .O(n211) );
  NR2T U1406 ( .I1(n2383), .I2(n282), .O(n1174) );
  ND3P U1407 ( .I1(n1044), .I2(n215), .I3(n1919), .O(n205) );
  AOI13HS U1408 ( .B1(n282), .B2(n1175), .B3(n831), .A1(n1176), .O(n1163) );
  MOAI1 U1409 ( .A1(n285), .A2(n2389), .B1(n2384), .B2(n1169), .O(n1175) );
  INV2 U1410 ( .I(n272), .O(n1176) );
  NR2T U1411 ( .I1(n590), .I2(n580), .O(n1024) );
  ND3 U1412 ( .I1(n548), .I2(n17), .I3(n1114), .O(n23) );
  OAI12 U1413 ( .B1(n1742), .B2(n1737), .A1(n1743), .O(n79) );
  ND3 U1414 ( .I1(n1744), .I2(n2377), .I3(n972), .O(n1743) );
  AOI12S U1415 ( .B1(n948), .B2(n2374), .A1(n1744), .O(n1742) );
  NR2 U1416 ( .I1(n2375), .I2(n709), .O(n705) );
  NR2T U1417 ( .I1(n2345), .I2(n605), .O(n614) );
  NR2T U1418 ( .I1(n2365), .I2(n2369), .O(n729) );
  NR2P U1419 ( .I1(n2276), .I2(n2281), .O(n659) );
  AOI13HS U1420 ( .B1(n896), .B2(n2334), .B3(n897), .A1(n898), .O(n893) );
  NR2 U1421 ( .I1(n536), .I2(n44), .O(n1542) );
  INV2 U1422 ( .I(n37), .O(n1541) );
  XNR2 U1423 ( .I1(n695), .I2(n101), .O(n1816) );
  NR2P U1424 ( .I1(n2322), .I2(n512), .O(n1274) );
  ND3P U1425 ( .I1(n809), .I2(n2392), .I3(n817), .O(n237) );
  OAI112 U1426 ( .C1(n389), .C2(n2267), .A1(n2268), .B1(n2269), .O(n1206) );
  OAI12S U1427 ( .B1(n1214), .B2(n1211), .A1(n2271), .O(n2268) );
  OR3B2 U1428 ( .I1(n2270), .B1(n380), .B2(n1213), .O(n2269) );
  ND3 U1429 ( .I1(n912), .I2(n918), .I3(n2082), .O(n1267) );
  NR2 U1430 ( .I1(n500), .I2(n2330), .O(n2082) );
  ND2P U1431 ( .I1(n1274), .I2(n2326), .O(n516) );
  ND3P U1432 ( .I1(n831), .I2(n2382), .I3(n840), .O(n265) );
  OAI12 U1433 ( .B1(n565), .B2(n14), .A1(n1106), .O(n19) );
  ND3 U1434 ( .I1(n18), .I2(n21), .I3(n1100), .O(n1106) );
  NR2P U1435 ( .I1(n2368), .I2(n958), .O(n706) );
  OAI12 U1436 ( .B1(n338), .B2(n2332), .A1(n335), .O(n340) );
  NR2P U1437 ( .I1(n122), .I2(n2430), .O(n139) );
  OA22 U1438 ( .A1(n374), .A2(n1218), .B1(n653), .B2(n387), .O(n1217) );
  AOI13HS U1439 ( .B1(n653), .B2(n656), .B3(n1208), .A1(n1219), .O(n1218) );
  NR3P U1440 ( .I1(n1220), .I2(n388), .I3(n659), .O(n1219) );
  XNR2 U1441 ( .I1(n653), .I2(n380), .O(n1220) );
  NR2 U1442 ( .I1(n2432), .I2(n2421), .O(n737) );
  ND3P U1443 ( .I1(n146), .I2(n2404), .I3(n793), .O(n165) );
  NR2P U1444 ( .I1(n774), .I2(n2413), .O(n162) );
  AOI13HS U1445 ( .B1(n2295), .B2(n1960), .B3(n657), .A1(n2296), .O(n2288) );
  INV2 U1446 ( .I(n659), .O(n2295) );
  NR3P U1447 ( .I1(n658), .I2(n1960), .I3(n2005), .O(n2296) );
  ND3 U1448 ( .I1(n605), .I2(n225), .I3(n1050), .O(n600) );
  ND3 U1449 ( .I1(n352), .I2(n1197), .I3(n2194), .O(n349) );
  INV2 U1450 ( .I(n254), .O(n817) );
  ND3 U1451 ( .I1(n2371), .I2(n62), .I3(n972), .O(n703) );
  NR2P U1452 ( .I1(n2350), .I2(n1016), .O(n1030) );
  NR2P U1453 ( .I1(n135), .I2(n2426), .O(n762) );
  NR2P U1454 ( .I1(n2416), .I2(n147), .O(n789) );
  BUF2 U1455 ( .I(n74), .O(n2379) );
  OAI12 U1458 ( .B1(n725), .B2(n726), .A1(n727), .O(n65) );
  INV2 U1459 ( .I(n729), .O(n726) );
  OAI112S U1460 ( .C1(n728), .C2(n706), .A1(n2365), .B1(n2379), .O(n727) );
  NR2 U1461 ( .I1(n2370), .I2(n709), .O(n728) );
  NR2P U1462 ( .I1(n474), .I2(n2320), .O(n2147) );
  ND3 U1463 ( .I1(n163), .I2(n2416), .I3(n448), .O(n456) );
  NR2P U1464 ( .I1(n2406), .I2(n774), .O(n1434) );
  ND3 U1465 ( .I1(n2364), .I2(n2357), .I3(n1004), .O(n669) );
  NR2P U1466 ( .I1(n2345), .I2(n1042), .O(n1055) );
  NR2P U1467 ( .I1(n2319), .I2(n471), .O(n2148) );
  ND3 U1468 ( .I1(n45), .I2(n1081), .I3(n1082), .O(n526) );
  BUF2 U1469 ( .I(n486), .O(n2318) );
  ND3 U1470 ( .I1(n551), .I2(n21), .I3(n1107), .O(n1492) );
  BUF2 U1471 ( .I(n421), .O(n2429) );
  ND3 U1472 ( .I1(n1110), .I2(n22), .I3(n1111), .O(n549) );
  BUF2 U1473 ( .I(n453), .O(n2412) );
  NR2 U1474 ( .I1(n1859), .I2(n192), .O(n1874) );
  ND3 U1475 ( .I1(n842), .I2(n2385), .I3(n1162), .O(n1156) );
  ND3 U1476 ( .I1(n840), .I2(n1161), .I3(n841), .O(n1157) );
  OA22 U1477 ( .A1(n834), .A2(n1159), .B1(n266), .B2(n1160), .O(n1158) );
  BUF2 U1478 ( .I(n123), .O(n2433) );
  AOI112P U1479 ( .C1(n860), .C2(n861), .A1(n307), .B1(n2338), .O(n859) );
  ND3 U1480 ( .I1(n862), .I2(n850), .I3(n2340), .O(n860) );
  ND3 U1481 ( .I1(n305), .I2(n304), .I3(n2344), .O(n861) );
  ND3 U1482 ( .I1(n382), .I2(n653), .I3(n650), .O(n379) );
  MOAI1P U1483 ( .A1(n615), .A2(n2348), .B1(n2348), .B2(n221), .O(n217) );
  BUF2 U1484 ( .I(n117), .O(n2423) );
  ND3 U1485 ( .I1(n1494), .I2(n1495), .I3(n1496), .O(n566) );
  ND3 U1486 ( .I1(n1111), .I2(n1095), .I3(n562), .O(n1494) );
  ND3 U1487 ( .I1(n548), .I2(n1102), .I3(n1105), .O(n1495) );
  OA22 U1488 ( .A1(n21), .A2(n1489), .B1(n557), .B2(n1492), .O(n1496) );
  ND3 U1489 ( .I1(n2341), .I2(n850), .I3(n865), .O(n864) );
  ND3 U1490 ( .I1(n2355), .I2(n996), .I3(n98), .O(n994) );
  ND3 U1491 ( .I1(n2417), .I2(n793), .I3(n794), .O(n151) );
  NR2 U1492 ( .I1(n2403), .I2(n2411), .O(n794) );
  OAI112S U1493 ( .C1(n918), .C2(n506), .A1(n516), .B1(n1273), .O(n1270) );
  ND2 U1494 ( .I1(n1274), .I2(n2324), .O(n1273) );
  BUF2 U1495 ( .I(n92), .O(n2360) );
  ND3 U1496 ( .I1(n338), .I2(n1329), .I3(n1330), .O(n1323) );
  OAI112S U1497 ( .C1(n961), .C2(n724), .A1(n962), .B1(n963), .O(n946) );
  ND3 U1498 ( .I1(n2369), .I2(n964), .I3(n71), .O(n962) );
  ND3 U1499 ( .I1(n1960), .I2(n2005), .I3(n374), .O(n2285) );
  ND3 U1500 ( .I1(n135), .I2(n736), .I3(n415), .O(n739) );
  INV2 U1501 ( .I(n1448), .O(n2469) );
  OAI112S U1502 ( .C1(n227), .C2(n1051), .A1(n1052), .B1(n1053), .O(n1046) );
  ND3 U1503 ( .I1(n605), .I2(n221), .I3(n204), .O(n1052) );
  AOI13HS U1504 ( .B1(n1054), .B2(n603), .B3(n1055), .A1(n1056), .O(n1053) );
  AOI112P U1505 ( .C1(n615), .C2(n1057), .A1(n204), .B1(n605), .O(n1056) );
  INV2 U1506 ( .I(n1446), .O(n2474) );
  OAI112S U1507 ( .C1(n1043), .C2(n1909), .A1(n1910), .B1(n1911), .O(n1908) );
  INV2 U1508 ( .I(n1055), .O(n1909) );
  ND3 U1509 ( .I1(n615), .I2(n2348), .I3(n222), .O(n1911) );
  ND3 U1510 ( .I1(n603), .I2(n221), .I3(n610), .O(n1910) );
  AOI112P U1511 ( .C1(n329), .C2(n330), .A1(n331), .B1(n332), .O(n327) );
  ND3 U1512 ( .I1(n77), .I2(n2366), .I3(n973), .O(n1752) );
  NR2P U1513 ( .I1(n605), .I2(n603), .O(n1919) );
  OAI12S U1514 ( .B1(n2358), .B2(n668), .A1(n669), .O(n667) );
  ND2 U1515 ( .I1(n1249), .I2(n468), .O(n1248) );
  ND3 U1516 ( .I1(n20), .I2(n2399), .I3(n1110), .O(n1489) );
  OAI12S U1517 ( .B1(n2371), .B2(n702), .A1(n703), .O(n701) );
  OAI12S U1518 ( .B1(n1670), .B2(n265), .A1(n273), .O(n1689) );
  OAI112S U1519 ( .C1(n2325), .C2(n516), .A1(n503), .B1(n1267), .O(n2081) );
  MOAI1 U1520 ( .A1(n43), .A2(n44), .B1(n45), .B2(n44), .O(n33) );
  ND2 U1521 ( .I1(n281), .I2(n1693), .O(n825) );
  ND3 U1522 ( .I1(n2385), .I2(n285), .I3(n1694), .O(n1693) );
  NR2 U1523 ( .I1(n2386), .I2(n282), .O(n1694) );
  INV2 U1524 ( .I(n2276), .O(n389) );
  NR2P U1525 ( .I1(n162), .I2(n793), .O(n452) );
  MOAI1 U1526 ( .A1(n20), .A2(n21), .B1(n22), .B2(n21), .O(n10) );
  AOI12S U1527 ( .B1(n2337), .B2(n1305), .A1(n315), .O(n1296) );
  ND3 U1528 ( .I1(n368), .I2(n1198), .I3(n627), .O(n1191) );
  AO222 U1529 ( .A1(n634), .A2(n1199), .B1(n1200), .B2(n361), .C1(n629), .C2(
        n632), .O(n1198) );
  NR2 U1530 ( .I1(n632), .I2(n366), .O(n1200) );
  OAI12S U1531 ( .B1(n352), .B2(n624), .A1(n1201), .O(n1199) );
  INV2 U1532 ( .I(n1448), .O(n2470) );
  INV2 U1533 ( .I(n1446), .O(n2475) );
  INV2 U1534 ( .I(n1381), .O(n2485) );
  INV2 U1535 ( .I(n1379), .O(n2491) );
  ND3 U1536 ( .I1(n1800), .I2(n2006), .I3(n659), .O(n387) );
  ND3 U1537 ( .I1(n806), .I2(n257), .I3(n1628), .O(n1627) );
  NR2 U1538 ( .I1(n254), .I2(n252), .O(n1628) );
  INV2 U1539 ( .I(n702), .O(n707) );
  ND3 U1540 ( .I1(n773), .I2(n2408), .I3(n2414), .O(n772) );
  MOAI1 U1541 ( .A1(n774), .A2(n442), .B1(n443), .B2(n2404), .O(n773) );
  ND3 U1542 ( .I1(n305), .I2(n306), .I3(n2342), .O(n298) );
  MOAI1 U1543 ( .A1(n307), .A2(n308), .B1(n309), .B2(n310), .O(n306) );
  OAI12S U1544 ( .B1(n2343), .B2(n312), .A1(n303), .O(n310) );
  OAI12S U1545 ( .B1(n119), .B2(n2430), .A1(n121), .O(n118) );
  OA12 U1546 ( .B1(n122), .B2(n2433), .A1(n124), .O(n119) );
  AOI12 U1547 ( .B1(n1087), .B2(n1546), .A1(n2394), .O(n1545) );
  ND2 U1548 ( .I1(n1071), .I2(n45), .O(n1546) );
  ND3 U1549 ( .I1(n2361), .I2(n2353), .I3(n1005), .O(n1814) );
  ND3 U1551 ( .I1(n2356), .I2(n680), .I3(n681), .O(n678) );
  NR2 U1553 ( .I1(n2363), .I2(n682), .O(n681) );
  AN3 U1554 ( .I1(n243), .I2(n1614), .I3(n1621), .O(n1141) );
  NR2 U1555 ( .I1(n2391), .I2(n252), .O(n1621) );
  AN3 U1556 ( .I1(n1670), .I2(n270), .I3(n1691), .O(n1168) );
  NR2 U1557 ( .I1(n2386), .I2(n2380), .O(n1691) );
  AN3 U1558 ( .I1(n1327), .I2(n338), .I3(n1328), .O(n328) );
  NR2 U1559 ( .I1(n323), .I2(n334), .O(n1328) );
  AN3 U1560 ( .I1(n382), .I2(n1800), .I3(n1212), .O(n651) );
  ND3 U1561 ( .I1(n713), .I2(n2376), .I3(n714), .O(n712) );
  NR2 U1562 ( .I1(n2370), .I2(n715), .O(n714) );
  AOI12S U1563 ( .B1(n1120), .B2(n1481), .A1(n2399), .O(n1480) );
  ND2 U1564 ( .I1(n1100), .I2(n2401), .O(n1481) );
  OAI12S U1565 ( .B1(n1275), .B2(n1276), .A1(n500), .O(n1268) );
  NR2 U1566 ( .I1(n2329), .I2(n1277), .O(n1275) );
  AOI13HS U1567 ( .B1(n511), .B2(n512), .B3(n919), .A1(n1278), .O(n1277) );
  NR2 U1568 ( .I1(n511), .I2(n517), .O(n1278) );
  OA12 U1569 ( .B1(n149), .B2(n2414), .A1(n151), .O(n148) );
  AOI12S U1570 ( .B1(n2415), .B2(n2409), .A1(n154), .O(n149) );
  NR2 U1571 ( .I1(n513), .I2(n2070), .O(n2077) );
  INV2 U1572 ( .I(n1082), .O(n1559) );
  INV2 U1573 ( .I(n1503), .O(n1442) );
  AN3 U1574 ( .I1(n129), .I2(n2429), .I3(n139), .O(n426) );
  INV2 U1575 ( .I(n1505), .O(n1444) );
  INV2 U1576 ( .I(n1111), .O(n1493) );
  ND3 U1577 ( .I1(n211), .I2(n216), .I3(n1913), .O(n1907) );
  ND3 U1578 ( .I1(n215), .I2(n225), .I3(n226), .O(n1913) );
  OA22 U1579 ( .A1(n274), .A2(n265), .B1(n275), .B2(n276), .O(n271) );
  ND2 U1580 ( .I1(n1186), .I2(n2200), .O(n353) );
  OA22 U1581 ( .A1(n1166), .A2(n282), .B1(n2385), .B2(n273), .O(n1165) );
  AOI12S U1582 ( .B1(n831), .B2(n1167), .A1(n1168), .O(n1166) );
  OAI12S U1583 ( .B1(n270), .B2(n1169), .A1(n267), .O(n1167) );
  INV2 U1584 ( .I(n1120), .O(n1114) );
  INV2 U1585 ( .I(n2070), .O(n2061) );
  OA22 U1586 ( .A1(n2408), .A2(n456), .B1(n147), .B2(n165), .O(n1433) );
  OA222 U1587 ( .A1(n276), .A2(n285), .B1(n274), .B2(n838), .C1(n282), .C2(
        n267), .O(n828) );
  INV2 U1588 ( .I(n1906), .O(n1051) );
  NR2 U1589 ( .I1(n215), .I2(n224), .O(n223) );
  OA22 U1590 ( .A1(n246), .A2(n237), .B1(n247), .B2(n248), .O(n242) );
  ND2 U1591 ( .I1(n1209), .I2(n2276), .O(n381) );
  ND2 U1592 ( .I1(n841), .I2(n842), .O(n283) );
  INV2 U1593 ( .I(n2024), .O(n883) );
  NR2 U1594 ( .I1(n1692), .I2(n2380), .O(n1690) );
  AOI13HS U1595 ( .B1(n834), .B2(n2387), .B3(n1174), .A1(n269), .O(n1692) );
  NR2 U1596 ( .I1(n1151), .I2(n1152), .O(n1150) );
  OAI112S U1597 ( .C1(n824), .C2(n1163), .A1(n1164), .B1(n1165), .O(n1151) );
  ND3 U1598 ( .I1(n278), .I2(n1153), .I3(n1154), .O(n1152) );
  ND3 U1599 ( .I1(n1170), .I2(n2388), .I3(n824), .O(n1164) );
  INV2 U1600 ( .I(n1050), .O(n1917) );
  NR2 U1601 ( .I1(n598), .I2(n599), .O(n597) );
  AOI13HS U1602 ( .B1(n600), .B2(n216), .B3(n601), .A1(n2346), .O(n598) );
  ND3 U1603 ( .I1(n603), .I2(n221), .I3(n604), .O(n601) );
  NR2 U1604 ( .I1(n605), .I2(n215), .O(n604) );
  ND2 U1605 ( .I1(n485), .I2(n2318), .O(n476) );
  OA12 U1606 ( .B1(n282), .B2(n833), .A1(n281), .O(n832) );
  OA12 U1607 ( .B1(n270), .B2(n834), .A1(n835), .O(n833) );
  ND3 U1608 ( .I1(n824), .I2(n2381), .I3(n270), .O(n835) );
  ND2 U1609 ( .I1(n224), .I2(n2347), .O(n1057) );
  NR2 U1610 ( .I1(n455), .I2(n2416), .O(n454) );
  INV2 U1611 ( .I(n157), .O(n156) );
  NR2 U1612 ( .I1(n129), .I2(n130), .O(n126) );
  INV2 U1613 ( .I(n128), .O(n127) );
  INV2 U1614 ( .I(n2327), .O(n508) );
  ND2 U1615 ( .I1(n2326), .I2(n2322), .O(n504) );
  BUF2 U1616 ( .I(n2516), .O(n2505) );
  BUF2 U1617 ( .I(n2516), .O(n2506) );
  BUF2 U1618 ( .I(n2514), .O(n2509) );
  BUF2 U1619 ( .I(n2514), .O(n2510) );
  ND3 U1620 ( .I1(n1221), .I2(n380), .I3(n1213), .O(n394) );
  BUF2 U1621 ( .I(n2515), .O(n2508) );
  BUF2 U1622 ( .I(n2513), .O(n2511) );
  ND2 U1623 ( .I1(n814), .I2(n806), .O(n807) );
  INV2 U1624 ( .I(n1381), .O(n2486) );
  NR2 U1625 ( .I1(n319), .I2(n338), .O(n1326) );
  BUF1 U1626 ( .I(n2539), .O(n2537) );
  BUF1 U1627 ( .I(n2539), .O(n2538) );
  BUF1 U1628 ( .I(n2539), .O(n2536) );
  BUF1 U1629 ( .I(n2513), .O(n2512) );
  INV3 U1630 ( .I(n2544), .O(n2541) );
  INV3 U1631 ( .I(n2543), .O(n2542) );
  INV3 U1632 ( .I(n2545), .O(n2540) );
  XOR2P U1633 ( .I1(n1992), .I2(n1780), .O(n862) );
  MOAI1 U1634 ( .A1(n2505), .A2(n1828), .B1(n1567), .B2(n2509), .O(n1992) );
  XOR2P U1635 ( .I1(n2256), .I2(n1898), .O(n366) );
  MOAI1 U1636 ( .A1(n2506), .A2(n1882), .B1(n1386), .B2(n2510), .O(n2256) );
  XOR2P U1637 ( .I1(n1996), .I2(n1997), .O(n1294) );
  MOAI1 U1638 ( .A1(n2501), .A2(n1842), .B1(n1998), .B2(n2502), .O(n1996) );
  BUF2 U1639 ( .I(n2169), .O(n2446) );
  BUF2 U1640 ( .I(n2169), .O(n2447) );
  BUF2 U1641 ( .I(n2170), .O(n2443) );
  AO2222 U1642 ( .A1(n2495), .A2(n1990), .B1(n2492), .B2(n1991), .C1(n2487), 
        .C2(n1995), .D1(n2482), .D2(n1843), .O(n1842) );
  ND2P U1643 ( .I1(decrypt_shift[0]), .I2(n2260), .O(n2171) );
  ND2P U1644 ( .I1(n2259), .I2(n2260), .O(n2172) );
  XOR2P U1645 ( .I1(n1838), .I2(n1780), .O(n674) );
  MOAI1 U1646 ( .A1(n1839), .A2(n2498), .B1(n1840), .B2(n2502), .O(n1838) );
  AO2222 U1647 ( .A1(n2495), .A2(n1574), .B1(n2492), .B2(n1575), .C1(n2487), 
        .C2(n1837), .D1(n2482), .D2(n1836), .O(n1840) );
  XOR2P U1648 ( .I1(n1779), .I2(n1780), .O(n709) );
  MOAI1 U1649 ( .A1(n1781), .A2(n2530), .B1(n1782), .B2(n2535), .O(n1779) );
  XOR2P U1650 ( .I1(n1889), .I2(n1395), .O(n1859) );
  AO22 U1651 ( .A1(n2511), .A2(n1662), .B1(n1638), .B2(n2504), .O(n1889) );
  XOR2P U1652 ( .I1(n1529), .I2(n1398), .O(n17) );
  MOAI1 U1653 ( .A1(n1530), .A2(n2530), .B1(n1531), .B2(n2535), .O(n1529) );
  AO2222 U1654 ( .A1(n2479), .A2(n1532), .B1(n2476), .B2(n1533), .C1(n2471), 
        .C2(n1534), .D1(n2466), .D2(n1535), .O(n1531) );
  XOR2P U1655 ( .I1(n1460), .I2(n1395), .O(n774) );
  MOAI1 U1656 ( .A1(n2518), .A2(n1439), .B1(n2528), .B2(n1461), .O(n1460) );
  AO2222 U1657 ( .A1(n2479), .A2(n1459), .B1(n2476), .B2(n1443), .C1(n2471), 
        .C2(n1445), .D1(n2466), .D2(n1447), .O(n1461) );
  XOR2P U1658 ( .I1(n1892), .I2(n1893), .O(n590) );
  MOAI1 U1660 ( .A1(n2505), .A2(n1650), .B1(n1883), .B2(n2509), .O(n1892) );
  XOR2P U1661 ( .I1(n2174), .I2(n1649), .O(n468) );
  MOAI1 U1662 ( .A1(n2507), .A2(n2000), .B1(n1570), .B2(n2508), .O(n2174) );
  XOR2P U1663 ( .I1(n2220), .I2(n1881), .O(n634) );
  AO22 U1664 ( .A1(n2504), .A2(n2221), .B1(n1626), .B2(n2512), .O(n2220) );
  XOR2P U1665 ( .I1(n2175), .I2(n1624), .O(n484) );
  MOAI1 U1666 ( .A1(n2507), .A2(n2176), .B1(n2177), .B2(n2509), .O(n2175) );
  XOR2P U1667 ( .I1(n1623), .I2(n1624), .O(n814) );
  MOAI1 U1668 ( .A1(n2499), .A2(n1625), .B1(n1626), .B2(n2503), .O(n1623) );
  MOAI1 U1669 ( .A1(n2500), .A2(n1885), .B1(n1404), .B2(n2501), .O(n1884) );
  NR3P U1670 ( .I1(n2397), .I2(n1083), .I3(n49), .O(n1073) );
  NR3P U1671 ( .I1(n603), .I2(n605), .I3(n1912), .O(n1918) );
  NR3P U1672 ( .I1(n691), .I2(n2362), .I3(n675), .O(n991) );
  NR3P U1673 ( .I1(n2401), .I2(n1112), .I3(n25), .O(n1102) );
  AOI112P U1674 ( .C1(n1066), .C2(n1067), .A1(n1068), .B1(n1069), .O(n543) );
  AO13 U1675 ( .B1(n2397), .B2(n1070), .B3(n1071), .A1(n1072), .O(n1069) );
  AO22 U1676 ( .A1(n538), .A2(n38), .B1(n2395), .B2(n1076), .O(n1070) );
  AN2 U1677 ( .I1(n1073), .I2(n1074), .O(n1072) );
  AOI112P U1678 ( .C1(n1095), .C2(n1096), .A1(n1097), .B1(n1098), .O(n567) );
  AO13 U1679 ( .B1(n2401), .B2(n1099), .B3(n1100), .A1(n1101), .O(n1098) );
  AO22 U1680 ( .A1(n562), .A2(n16), .B1(n2399), .B2(n1105), .O(n1099) );
  AN2 U1681 ( .I1(n1102), .I2(n1103), .O(n1101) );
  MOAI1 U1682 ( .A1(n2500), .A2(n1650), .B1(n1400), .B2(n2502), .O(n1648) );
  MOAI1 U1683 ( .A1(n2501), .A2(n1580), .B1(n2003), .B2(n2502), .O(n2168) );
  INV3 U1684 ( .I(n502), .O(n513) );
  MOAI1 U1685 ( .A1(n2506), .A2(n1570), .B1(n2511), .B2(n1571), .O(n1569) );
  AO2222 U1686 ( .A1(n2496), .A2(n1572), .B1(n2493), .B2(n1573), .C1(n2488), 
        .C2(n1574), .D1(n2483), .D2(n1575), .O(n1571) );
  XNR2 U1687 ( .I1(n1661), .I2(n1722), .O(n1720) );
  XNR2 U1688 ( .I1(n1661), .I2(n1662), .O(n1659) );
  INV3 U1689 ( .I(n877), .O(n338) );
  INV3 U1690 ( .I(n890), .O(n332) );
  MOAI1 U1691 ( .A1(n2506), .A2(n1989), .B1(n1998), .B2(n2510), .O(n2173) );
  MOAI1 U1692 ( .A1(n2519), .A2(n1501), .B1(n2528), .B2(n1502), .O(n1500) );
  MOAI1 U1693 ( .A1(n2499), .A2(n1385), .B1(n1386), .B2(n2503), .O(n1383) );
  INV3 U1694 ( .I(n1547), .O(n45) );
  MOAI1 U1695 ( .A1(n2499), .A2(n1403), .B1(n1631), .B2(n2503), .O(n1629) );
  ND3P U1696 ( .I1(n334), .I2(n877), .I3(n319), .O(n1317) );
  XOR2 U1697 ( .I1(n2257), .I2(n1637), .O(n369) );
  MOAI1 U1698 ( .A1(n2505), .A2(n1385), .B1(n1399), .B2(n2510), .O(n2257) );
  XOR2 U1699 ( .I1(n1401), .I2(n1402), .O(n427) );
  MOAI1 U1700 ( .A1(n2516), .A2(n1403), .B1(n1404), .B2(n2510), .O(n1401) );
  AOI22 U1701 ( .A1(n2504), .A2(n2177), .B1(n1825), .B2(n2512), .O(n1507) );
  MOAI1 U1702 ( .A1(n2500), .A2(n1583), .B1(n1577), .B2(n2502), .O(n1993) );
  INV3 U1703 ( .I(n499), .O(n500) );
  INV3 U1704 ( .I(n916), .O(n512) );
  NR2T U1705 ( .I1(n17), .I2(n25), .O(n1100) );
  NR2T U1706 ( .I1(n40), .I2(n49), .O(n1071) );
  NR2T U1707 ( .I1(n2394), .I2(n1547), .O(n538) );
  NR2T U1708 ( .I1(n674), .I2(n1002), .O(n1004) );
  NR2T U1709 ( .I1(n709), .I2(n970), .O(n972) );
  OR2 U1710 ( .I1(n1509), .I2(n1585), .O(n2004) );
  AO112 U1711 ( .C1(n2016), .C2(n877), .A1(n1312), .B1(n879), .O(n1509) );
  AO112 U1712 ( .C1(n334), .C2(n2007), .A1(n2008), .B1(n898), .O(n1585) );
  NR2T U1713 ( .I1(n2398), .I2(n1119), .O(n562) );
  ND3P U1714 ( .I1(n2362), .I2(n1002), .I3(n2364), .O(n668) );
  ND3P U1715 ( .I1(n77), .I2(n970), .I3(n62), .O(n702) );
  NR2T U1716 ( .I1(n337), .I2(n332), .O(n882) );
  NR2T U1717 ( .I1(n285), .I2(n837), .O(n1670) );
  OAI112 U1718 ( .C1(n1258), .C2(n2322), .A1(n1259), .B1(n1260), .O(n493) );
  ND2 U1719 ( .I1(n1261), .I2(n1262), .O(n1259) );
  AOI13HS U1720 ( .B1(n502), .B2(n2327), .B3(n1263), .A1(n1264), .O(n1258) );
  AOI112P U1721 ( .C1(n1265), .C2(n1266), .A1(n2326), .B1(n502), .O(n1264) );
  XOR2 U1722 ( .I1(n1454), .I2(n1388), .O(n453) );
  MOAI1 U1723 ( .A1(n2517), .A2(n1455), .B1(n2529), .B2(n1456), .O(n1454) );
  AO2222 U1724 ( .A1(n2479), .A2(n1457), .B1(n2476), .B2(n1458), .C1(n2471), 
        .C2(n1459), .D1(n2466), .D2(n1443), .O(n1456) );
  XOR2 U1726 ( .I1(n1387), .I2(n1388), .O(n421) );
  MOAI1 U1727 ( .A1(n2505), .A2(n1389), .B1(n2511), .B2(n1390), .O(n1387) );
  AO2222 U1728 ( .A1(n2496), .A2(n1391), .B1(n2493), .B2(n1392), .C1(n2488), 
        .C2(n1393), .D1(n2483), .D2(n1376), .O(n1390) );
  XOR2 U1729 ( .I1(n1827), .I2(n1769), .O(n92) );
  MOAI1 U1730 ( .A1(n2499), .A2(n1828), .B1(n1818), .B2(n2502), .O(n1827) );
  XOR2 U1731 ( .I1(n1880), .I2(n1881), .O(n192) );
  MOAI1 U1732 ( .A1(n2500), .A2(n1882), .B1(n1883), .B2(n2501), .O(n1880) );
  XOR2 U1733 ( .I1(n1988), .I2(n1514), .O(n863) );
  MOAI1 U1734 ( .A1(n2500), .A2(n1989), .B1(n1584), .B2(n2501), .O(n1988) );
  XOR2 U1735 ( .I1(n2178), .I2(n1769), .O(n486) );
  MOAI1 U1736 ( .A1(n2501), .A2(n2176), .B1(n1587), .B2(n2503), .O(n2178) );
  AOI13HS U1737 ( .B1(n417), .B2(n2420), .B3(n1367), .A1(n1368), .O(n1365) );
  AOI112P U1738 ( .C1(n1369), .C2(n1370), .A1(n135), .B1(n116), .O(n1368) );
  ND2 U1739 ( .I1(n758), .I2(n760), .O(n1369) );
  ND3 U1740 ( .I1(n130), .I2(n424), .I3(n409), .O(n1370) );
  XOR2 U1741 ( .I1(n2252), .I2(n2253), .O(n348) );
  AO22 U1742 ( .A1(n2511), .A2(n1389), .B1(n1900), .B2(n2504), .O(n2252) );
  XOR2 U1743 ( .I1(n1397), .I2(n1398), .O(n117) );
  AO22 U1744 ( .A1(n2504), .A2(n1399), .B1(n1400), .B2(n2512), .O(n1397) );
  OAI112 U1745 ( .C1(n2329), .C2(n2074), .A1(n2075), .B1(n2076), .O(n920) );
  ND3 U1746 ( .I1(n2067), .I2(n2066), .I3(n912), .O(n2076) );
  ND3 U1747 ( .I1(n2329), .I2(n513), .I3(n2061), .O(n2075) );
  AOI13HS U1748 ( .B1(n916), .B2(n2325), .B3(n1261), .A1(n2077), .O(n2074) );
  OA12 U1749 ( .B1(n99), .B2(n1813), .A1(n2354), .O(n1812) );
  AOI12S U1750 ( .B1(n2355), .B2(n682), .A1(n675), .O(n1813) );
  NR2T U1751 ( .I1(n378), .I2(n382), .O(n1213) );
  NR2T U1752 ( .I1(n354), .I2(n361), .O(n2194) );
  INV2 U1753 ( .I(n49), .O(n539) );
  ND3P U1754 ( .I1(n319), .I2(n894), .I3(n338), .O(n2021) );
  AOI112P U1755 ( .C1(n1114), .C2(n1112), .A1(n1115), .B1(n1116), .O(n1113) );
  INV2 U1756 ( .I(n23), .O(n1116) );
  AOI13HS U1757 ( .B1(n1117), .B2(n560), .B3(n1118), .A1(n1119), .O(n1115) );
  OAI112S U1758 ( .C1(n1095), .C2(n1100), .A1(n2398), .B1(n2401), .O(n1117) );
  AOI112P U1759 ( .C1(n685), .C2(n93), .A1(n686), .B1(n687), .O(n684) );
  NR2 U1760 ( .I1(n675), .I2(n95), .O(n687) );
  NR2P U1761 ( .I1(n1547), .I2(n46), .O(n43) );
  ND2P U1762 ( .I1(decrypt_shift[3]), .I2(decrypt_shift[2]), .O(n1640) );
  OA112 U1763 ( .C1(n2063), .C2(n2328), .A1(n2064), .B1(n2065), .O(n1260) );
  ND3 U1764 ( .I1(n2066), .I2(n2323), .I3(n1263), .O(n2065) );
  ND3 U1765 ( .I1(n2067), .I2(n513), .I3(n1262), .O(n2064) );
  AOI13HS U1766 ( .B1(n2067), .B2(n502), .B3(n912), .A1(n2068), .O(n2063) );
  BUF2 U1767 ( .I(n679), .O(n2355) );
  BUF2 U1768 ( .I(n1075), .O(n2394) );
  AO2222 U1769 ( .A1(n2495), .A2(n1831), .B1(n2492), .B2(n1819), .C1(n2487), 
        .C2(n1820), .D1(n2482), .D2(n1821), .O(n1828) );
  AO2222 U1770 ( .A1(n2495), .A2(n1654), .B1(n2492), .B2(n1895), .C1(n2487), 
        .C2(n1896), .D1(n2482), .D2(n1894), .O(n1650) );
  AO2222 U1771 ( .A1(n2495), .A2(n1633), .B1(n2492), .B2(n1634), .C1(n2487), 
        .C2(n1635), .D1(n2482), .D2(n1886), .O(n1625) );
  AO2222 U1772 ( .A1(n2495), .A2(n1995), .B1(n2492), .B2(n1843), .C1(n2487), 
        .C2(n1844), .D1(n2482), .D2(n1845), .O(n1583) );
  AO2222 U1773 ( .A1(n2495), .A2(n1653), .B1(n2492), .B2(n1654), .C1(n2487), 
        .C2(n1895), .D1(n2482), .D2(n1896), .O(n1882) );
  AO2222 U1774 ( .A1(n2496), .A2(n1632), .B1(n2493), .B2(n1633), .C1(n2488), 
        .C2(n1634), .D1(n2483), .D2(n1635), .O(n1403) );
  AO2222 U1775 ( .A1(n2495), .A2(n1991), .B1(n2492), .B2(n1995), .C1(n2487), 
        .C2(n1843), .D1(n2482), .D2(n1844), .O(n1989) );
  AO2222 U1776 ( .A1(n2495), .A2(n1829), .B1(n2492), .B2(n1830), .C1(n2487), 
        .C2(n1831), .D1(n2482), .D2(n1819), .O(n1580) );
  AO2222 U1777 ( .A1(n2495), .A2(n1652), .B1(n2492), .B2(n1653), .C1(n2487), 
        .C2(n1654), .D1(n2482), .D2(n1895), .O(n1385) );
  AO2222 U1778 ( .A1(n2495), .A2(n1888), .B1(n2492), .B2(n1632), .C1(n2487), 
        .C2(n1633), .D1(n2482), .D2(n1634), .O(n1885) );
  NR2P U1779 ( .I1(n890), .I2(n337), .O(n341) );
  AO2222 U1780 ( .A1(n2495), .A2(n2180), .B1(n2492), .B2(n1591), .C1(n2487), 
        .C2(n1590), .D1(n2482), .D2(n1589), .O(n2176) );
  AO2222 U1781 ( .A1(n2495), .A2(n1573), .B1(n2492), .B2(n1574), .C1(n2487), 
        .C2(n1575), .D1(n2482), .D2(n1837), .O(n2000) );
  BUF2 U1782 ( .I(n679), .O(n2356) );
  NR2P U1783 ( .I1(n613), .I2(n1054), .O(n1906) );
  ND2P U1784 ( .I1(decrypt_shift[3]), .I2(n2258), .O(n1642) );
  INV2 U1785 ( .I(n354), .O(n627) );
  INV2 U1786 ( .I(n378), .O(n648) );
  BUF2 U1787 ( .I(n723), .O(n2369) );
  BUF2 U1788 ( .I(n723), .O(n2368) );
  INV2 U1789 ( .I(n40), .O(n1083) );
  NR2P U1790 ( .I1(n424), .I2(n2424), .O(n758) );
  AO2222 U1791 ( .A1(n2495), .A2(n1830), .B1(n2492), .B2(n1831), .C1(n2487), 
        .C2(n1819), .D1(n2482), .D2(n1820), .O(n1568) );
  BUF2 U1792 ( .I(n2170), .O(n2442) );
  ND3P U1797 ( .I1(n2346), .I2(n214), .I3(n1906), .O(n1045) );
  BUF2 U1803 ( .I(n85), .O(n2354) );
  NR2P U1804 ( .I1(n655), .I2(n648), .O(n1208) );
  NR2P U1805 ( .I1(n2258), .I2(decrypt_shift[3]), .O(n1379) );
  NR2P U1806 ( .I1(n335), .I2(n894), .O(n2029) );
  BUF2 U1807 ( .I(n2169), .O(n2448) );
  NR2P U1808 ( .I1(n890), .I2(n897), .O(n1327) );
  BUF2 U1809 ( .I(n2170), .O(n2444) );
  ND3 U1810 ( .I1(n509), .I2(n916), .I3(n2330), .O(n497) );
  AO12 U1811 ( .B1(n1644), .B2(n980), .A1(n1646), .O(n88) );
  OAI22 U1812 ( .A1(n993), .A2(n102), .B1(n990), .B2(n668), .O(n1644) );
  AN3 U1813 ( .I1(n989), .I2(n675), .I3(n985), .O(n1646) );
  MOAI1P U1814 ( .A1(n1923), .A2(n615), .B1(n1924), .B2(n1925), .O(n599) );
  OAI12S U1815 ( .B1(n215), .B2(n228), .A1(n1926), .O(n1925) );
  OA13 U1816 ( .B1(n1043), .B2(n204), .B3(n214), .A1(n1914), .O(n1923) );
  ND3 U1817 ( .I1(n215), .I2(n613), .I3(n1054), .O(n1926) );
  NR2 U1818 ( .I1(n346), .I2(n347), .O(n345) );
  OAI112S U1819 ( .C1(n2314), .C2(n349), .A1(n350), .B1(n351), .O(n347) );
  AOI13HS U1820 ( .B1(n357), .B2(n360), .B3(n361), .A1(n362), .O(n358) );
  BUF2 U1821 ( .I(n458), .O(n2404) );
  BUF2 U1822 ( .I(n152), .O(n2415) );
  BUF2 U1823 ( .I(n579), .O(n2350) );
  BUF2 U1824 ( .I(n602), .O(n2345) );
  OA12 U1825 ( .B1(n1348), .B2(n130), .A1(n1349), .O(n748) );
  ND3 U1826 ( .I1(n1350), .I2(n424), .I3(n1351), .O(n1349) );
  AOI13HS U1827 ( .B1(n2427), .B2(n2423), .B3(n1352), .A1(n1353), .O(n1348) );
  XNR2 U1828 ( .I1(n2427), .I2(n2429), .O(n1350) );
  AO2222 U1829 ( .A1(n2495), .A2(n1843), .B1(n2492), .B2(n1844), .C1(n2487), 
        .C2(n1845), .D1(n2482), .D2(n1846), .O(n1578) );
  BUF2 U1830 ( .I(n496), .O(n2325) );
  MOAI1 U1831 ( .A1(n36), .A2(n37), .B1(n38), .B2(n39), .O(n34) );
  AO12 U1832 ( .B1(n40), .B2(n41), .A1(n42), .O(n39) );
  BUF2 U1833 ( .I(n836), .O(n2382) );
  ND3 U1834 ( .I1(n695), .I2(n675), .I3(n1798), .O(n1796) );
  OA112 U1835 ( .C1(n215), .C2(n1037), .A1(n1038), .B1(n1039), .O(n606) );
  OR3B2 U1836 ( .I1(n1043), .B1(n1044), .B2(n614), .O(n1038) );
  OA22 U1837 ( .A1(n613), .A2(n1040), .B1(n2349), .B2(n1045), .O(n1037) );
  OR3 U1838 ( .I1(n1040), .I2(n1041), .I3(n1042), .O(n1039) );
  BUF2 U1839 ( .I(n2169), .O(n2449) );
  BUF2 U1840 ( .I(n2170), .O(n2445) );
  BUF1 U1841 ( .I(n390), .O(n1801) );
  ND3 U1842 ( .I1(n1537), .I2(n523), .I3(n1538), .O(n1536) );
  NR2 U1843 ( .I1(n1068), .I2(n50), .O(n1537) );
  OA222 U1844 ( .A1(n48), .A2(n539), .B1(n1539), .B2(n38), .C1(n1540), .C2(n46), .O(n1538) );
  AOI13S U1845 ( .B1(n40), .B2(n1544), .B3(n2395), .A1(n1545), .O(n1539) );
  ND3 U1846 ( .I1(n1664), .I2(n1665), .I3(n1666), .O(n1663) );
  MAOI1 U1847 ( .A1(n837), .A2(n825), .B1(n831), .B2(n839), .O(n1664) );
  AOI112P U1848 ( .C1(n1689), .C2(n2384), .A1(n1690), .B1(n1168), .O(n1665) );
  AOI112P U1849 ( .C1(n286), .C2(n285), .A1(n826), .B1(n1155), .O(n1666) );
  ND3 U1850 ( .I1(n873), .I2(n874), .I3(n875), .O(n872) );
  AOI13HS U1851 ( .B1(n885), .B2(n337), .B3(n319), .A1(n886), .O(n874) );
  OA22 U1852 ( .A1(n893), .A2(n894), .B1(n2335), .B2(n895), .O(n873) );
  OA112 U1853 ( .C1(n876), .C2(n877), .A1(n878), .B1(n322), .O(n875) );
  INV2 U1854 ( .I(decrypt_shift[0]), .O(n2259) );
  INV2 U1855 ( .I(decrypt_shift[2]), .O(n2258) );
  XOR2P U1856 ( .I1(n1394), .I2(n1395), .O(n122) );
  MOAI1 U1857 ( .A1(n2509), .A2(n1372), .B1(n2511), .B2(n1396), .O(n1394) );
  AO2222 U1858 ( .A1(n2496), .A2(n1393), .B1(n2493), .B2(n1376), .C1(n2488), 
        .C2(n1378), .D1(n2483), .D2(n1380), .O(n1396) );
  XOR2P U1859 ( .I1(n1897), .I2(n1898), .O(n580) );
  MOAI1 U1860 ( .A1(n2506), .A2(n1625), .B1(n1631), .B2(n2509), .O(n1897) );
  BUF1 U1861 ( .I(n377), .O(n1817) );
  ND3 U1862 ( .I1(n2262), .I2(n2263), .I3(n2264), .O(n2261) );
  OA22 U1863 ( .A1(n1225), .A2(n2293), .B1(n1801), .B2(n381), .O(n2262) );
  OA222 U1864 ( .A1(n374), .A2(n2288), .B1(n386), .B2(n2289), .C1(n648), .C2(
        n2290), .O(n2263) );
  AOI112P U1865 ( .C1(n2265), .C2(n2005), .A1(n2266), .B1(n1206), .O(n2264) );
  BUF1 U1866 ( .I(n1104), .O(n2398) );
  ND2 U1867 ( .I1(n1686), .I2(n1687), .O(n286) );
  ND3 U1868 ( .I1(n824), .I2(n2381), .I3(n1674), .O(n1687) );
  ND3 U1869 ( .I1(n1688), .I2(n837), .I3(n270), .O(n1686) );
  MOAI1 U1870 ( .A1(n2000), .A2(n2498), .B1(n2504), .B2(n1839), .O(n1999) );
  INV2 U1871 ( .I(n970), .O(n74) );
  MOAI1 U1872 ( .A1(n2506), .A2(n1885), .B1(n2221), .B2(n2509), .O(n2254) );
  MOAI1 U1873 ( .A1(n2506), .A2(n1568), .B1(n2003), .B2(n2509), .O(n2001) );
  AN3 U1874 ( .I1(n1929), .I2(n1930), .I3(n1931), .O(n607) );
  ND3 U1875 ( .I1(n612), .I2(n1042), .I3(n614), .O(n1930) );
  OR3B2 U1876 ( .I1(n1045), .B1(n2348), .B2(n1041), .O(n1929) );
  AOI13HS U1877 ( .B1(n1924), .B2(n1912), .B3(n1050), .A1(n1932), .O(n1931) );
  OAI12S U1878 ( .B1(n2215), .B2(n362), .A1(n2313), .O(n2212) );
  AN2 U1879 ( .I1(n354), .I2(n628), .O(n2215) );
  OR3B2 U1880 ( .I1(n493), .B1(n494), .B2(n495), .O(n492) );
  OA222 U1881 ( .A1(n2324), .A2(n497), .B1(n498), .B2(n499), .C1(n500), .C2(
        n501), .O(n495) );
  OA222 U1882 ( .A1(n513), .A2(n516), .B1(n512), .B2(n517), .C1(n506), .C2(
        n518), .O(n498) );
  OA222 U1883 ( .A1(n502), .A2(n503), .B1(n504), .B2(n505), .C1(n506), .C2(
        n507), .O(n501) );
  ND2 U1884 ( .I1(n912), .I2(n499), .O(n1266) );
  INV2 U1885 ( .I(n167), .O(n150) );
  OA222 U1886 ( .A1(n45), .A2(n536), .B1(n537), .B2(n2397), .C1(n538), .C2(n37), .O(n527) );
  AOI112P U1887 ( .C1(n539), .C2(n41), .A1(n32), .B1(n540), .O(n537) );
  NR2 U1888 ( .I1(n40), .I2(n541), .O(n540) );
  ND3 U1889 ( .I1(n902), .I2(n903), .I3(n904), .O(n901) );
  NR2 U1890 ( .I1(n920), .I2(n493), .O(n902) );
  OA222 U1891 ( .A1(n905), .A2(n499), .B1(n906), .B2(n2326), .C1(n500), .C2(
        n907), .O(n904) );
  OA13 U1892 ( .B1(n908), .B2(n500), .B3(n909), .A1(n910), .O(n906) );
  BUF1 U1893 ( .I(n1320), .O(n2333) );
  NR2 U1894 ( .I1(n1203), .I2(n1204), .O(n1202) );
  ND3 U1895 ( .I1(n1215), .I2(n1216), .I3(n1217), .O(n1203) );
  OR3B2 U1896 ( .I1(n1205), .B1(n396), .B2(n643), .O(n1204) );
  OR3B2 U1897 ( .I1(n383), .B1(n1221), .B2(n655), .O(n1216) );
  NR2 U1898 ( .I1(n2057), .I2(n2058), .O(n2056) );
  AO222 U1899 ( .A1(n513), .A2(n2079), .B1(n2080), .B2(n2327), .C1(n2081), 
        .C2(n502), .O(n2057) );
  ND3 U1900 ( .I1(n494), .I2(n1260), .I3(n903), .O(n2058) );
  OAI12S U1901 ( .B1(n499), .B2(n909), .A1(n910), .O(n2080) );
  NR2 U1902 ( .I1(n1336), .I2(n1337), .O(n1335) );
  OAI112S U1903 ( .C1(n1364), .C2(n424), .A1(n1365), .B1(n1366), .O(n1336) );
  OAI112S U1904 ( .C1(n420), .C2(n124), .A1(n1338), .B1(n1339), .O(n1337) );
  OA22 U1905 ( .A1(n2423), .A2(n425), .B1(n2425), .B2(n137), .O(n1366) );
  NR2 U1906 ( .I1(n1034), .I2(n1035), .O(n1033) );
  AO2222 U1907 ( .A1(n1046), .A2(n1041), .B1(n1047), .B2(n2346), .C1(n226), 
        .C2(n612), .D1(n215), .D2(n1048), .O(n1034) );
  OAI112S U1908 ( .C1(n2346), .C2(n211), .A1(n606), .B1(n1036), .O(n1035) );
  INV2 U1909 ( .I(n600), .O(n1047) );
  ND3 U1910 ( .I1(n522), .I2(n523), .I3(n524), .O(n521) );
  OA222 U1911 ( .A1(n525), .A2(n526), .B1(n527), .B2(n38), .C1(n528), .C2(n46), 
        .O(n524) );
  NR2 U1912 ( .I1(n542), .I2(n51), .O(n522) );
  AOI112P U1913 ( .C1(n2396), .C2(n530), .A1(n35), .B1(n531), .O(n528) );
  ND3 U1914 ( .I1(n545), .I2(n546), .I3(n547), .O(n544) );
  OA222 U1915 ( .A1(n548), .A2(n549), .B1(n550), .B2(n16), .C1(n551), .C2(n552), .O(n547) );
  NR2 U1916 ( .I1(n566), .I2(n27), .O(n545) );
  AOI112P U1917 ( .C1(n2402), .C2(n554), .A1(n12), .B1(n555), .O(n552) );
  NR2 U1918 ( .I1(n423), .I2(n424), .O(n422) );
  ND3 U1919 ( .I1(n6), .I2(n7), .I3(n8), .O(n5) );
  OA22 U1920 ( .A1(n16), .A2(n23), .B1(n24), .B2(n25), .O(n7) );
  AOI112P U1921 ( .C1(n9), .C2(n10), .A1(n11), .B1(n12), .O(n8) );
  NR2 U1922 ( .I1(n26), .I2(n27), .O(n6) );
  ND3 U1923 ( .I1(n29), .I2(n30), .I3(n31), .O(n28) );
  MAOI1 U1924 ( .A1(n46), .A2(n47), .B1(n48), .B2(n49), .O(n30) );
  AOI112P U1925 ( .C1(n32), .C2(n33), .A1(n34), .B1(n35), .O(n31) );
  NR2 U1926 ( .I1(n50), .I2(n51), .O(n29) );
  NR2 U1927 ( .I1(n1254), .I2(n1255), .O(n1253) );
  OAI112S U1928 ( .C1(n502), .C2(n1267), .A1(n1268), .B1(n1269), .O(n1254) );
  OR3 U1929 ( .I1(n1256), .I2(n493), .I3(n1257), .O(n1255) );
  AOI13HS U1930 ( .B1(n502), .B2(n499), .B3(n1270), .A1(n1271), .O(n1269) );
  ND3 U1931 ( .I1(n1473), .I2(n546), .I3(n1474), .O(n1472) );
  OA222 U1932 ( .A1(n563), .A2(n24), .B1(n1475), .B2(n16), .C1(n551), .C2(
        n1476), .O(n1474) );
  NR2 U1933 ( .I1(n1097), .I2(n26), .O(n1473) );
  AOI13HS U1934 ( .B1(n1479), .B2(n2399), .B3(n17), .A1(n1480), .O(n1475) );
  INV1 U1935 ( .I(n675), .O(n90) );
  INV2 U1936 ( .I(n424), .O(n123) );
  ND2 U1937 ( .I1(n372), .I2(n373), .O(n371) );
  OA2222S U1938 ( .A1(n374), .A2(n375), .B1(n376), .B2(n1817), .C1(n378), .C2(
        n379), .D1(n380), .D2(n381), .O(n373) );
  OA112 U1939 ( .C1(n394), .C2(n2006), .A1(n395), .B1(n396), .O(n372) );
  AOI13HS U1940 ( .B1(n391), .B2(n1817), .B3(n382), .A1(n392), .O(n375) );
  AN3 U1941 ( .I1(n1918), .I2(n613), .I3(n610), .O(n1932) );
  ND2 U1942 ( .I1(n141), .I2(n142), .O(n140) );
  OA222 U1943 ( .A1(n143), .A2(n2407), .B1(n145), .B2(n146), .C1(n147), .C2(
        n148), .O(n142) );
  AOI112P U1944 ( .C1(n166), .C2(n167), .A1(n168), .B1(n169), .O(n141) );
  AOI13HS U1945 ( .B1(n2410), .B2(n2414), .B3(n155), .A1(n156), .O(n145) );
  AN2 U1946 ( .I1(n1548), .I2(n1549), .O(n48) );
  ND3 U1947 ( .I1(n1083), .I2(n1082), .I3(n1078), .O(n1548) );
  NR2 U1948 ( .I1(n2396), .I2(n46), .O(n1550) );
  AN2 U1949 ( .I1(n1482), .I2(n1483), .O(n24) );
  ND3 U1950 ( .I1(n1112), .I2(n1111), .I3(n1107), .O(n1482) );
  OR3B2 U1951 ( .I1(n556), .B1(n16), .B2(n1484), .O(n1483) );
  NR2 U1952 ( .I1(n1112), .I2(n2402), .O(n1484) );
  AN2 U1953 ( .I1(n167), .I2(n443), .O(n1430) );
  MOAI1 U1954 ( .A1(n1638), .A2(n2498), .B1(n1639), .B2(n2503), .O(n1636) );
  MOAI1 U1955 ( .A1(n1703), .A2(n2530), .B1(n1704), .B2(n2535), .O(n1702) );
  NR3P U1956 ( .I1(n335), .I2(n890), .I3(n331), .O(n898) );
  NR2T U1957 ( .I1(n44), .I2(n38), .O(n1082) );
  ND3P U1958 ( .I1(n44), .I2(n49), .I3(n1547), .O(n1087) );
  ND3P U1959 ( .I1(n512), .I2(n499), .I3(n2078), .O(n2070) );
  NR2 U1960 ( .I1(n2325), .I2(n2322), .O(n2078) );
  NR2T U1961 ( .I1(n16), .I2(n21), .O(n1111) );
  AOI13HS U1962 ( .B1(n2335), .B2(n890), .B3(n319), .A1(n2015), .O(n2014) );
  NR2 U1963 ( .I1(n890), .I2(n2334), .O(n2015) );
  ND2T U1964 ( .I1(encrypt_shift[3]), .I2(encrypt_shift[2]), .O(n1503) );
  AOI112P U1965 ( .C1(n1000), .C2(n1001), .A1(n2360), .B1(n990), .O(n999) );
  ND3 U1966 ( .I1(n675), .I2(n1002), .I3(n2357), .O(n1000) );
  ND2 U1967 ( .I1(n980), .I2(n2363), .O(n1001) );
  AOI112P U1968 ( .C1(n968), .C2(n969), .A1(n2374), .B1(n958), .O(n967) );
  ND3 U1969 ( .I1(n970), .I2(n2377), .I3(n2371), .O(n968) );
  ND2 U1970 ( .I1(n948), .I2(n2379), .O(n969) );
  AOI13HS U1971 ( .B1(n2410), .B2(n163), .B3(n439), .A1(n440), .O(n438) );
  NR2 U1972 ( .I1(n441), .I2(n442), .O(n440) );
  AOI112P U1973 ( .C1(n1436), .C2(n1437), .A1(n167), .B1(n146), .O(n1435) );
  ND2 U1974 ( .I1(n789), .I2(n791), .O(n1436) );
  ND3 U1975 ( .I1(n158), .I2(n2415), .I3(n441), .O(n1437) );
  AOI112P U1976 ( .C1(n887), .C2(n888), .A1(n319), .B1(n334), .O(n886) );
  ND3 U1977 ( .I1(n2336), .I2(n890), .I3(n877), .O(n887) );
  ND3 U1978 ( .I1(n332), .I2(n331), .I3(n338), .O(n888) );
  OAI12 U1979 ( .B1(n1804), .B2(n1799), .A1(n1805), .O(n106) );
  ND3 U1980 ( .I1(n1806), .I2(n675), .I3(n1004), .O(n1805) );
  AOI12S U1981 ( .B1(n980), .B2(n2359), .A1(n1806), .O(n1804) );
  ND2T U1982 ( .I1(encrypt_shift[3]), .I2(n2310), .O(n1505) );
  NR2 U1983 ( .I1(n674), .I2(n675), .O(n671) );
  ND3P U1984 ( .I1(n378), .I2(n2006), .I3(n380), .O(n383) );
  AOI112P U1985 ( .C1(n499), .C2(n1272), .A1(n909), .B1(n2328), .O(n1271) );
  ND2 U1986 ( .I1(n918), .I2(n513), .O(n1272) );
  AOI112P U1987 ( .C1(n45), .C2(n1085), .A1(n47), .B1(n1086), .O(n1084) );
  NR2 U1988 ( .I1(n40), .I2(n1087), .O(n1086) );
  OAI112S U1989 ( .C1(n2394), .C2(n37), .A1(n1088), .B1(n536), .O(n1085) );
  OAI112S U1990 ( .C1(n1066), .C2(n1071), .A1(n2394), .B1(n2396), .O(n1088) );
  ND3P U1991 ( .I1(n2315), .I2(n354), .I3(n352), .O(n363) );
  NR2T U1992 ( .I1(n1912), .I2(n1043), .O(n612) );
  BUF2 U1993 ( .I(n85), .O(n2353) );
  NR2P U1994 ( .I1(n502), .I2(n2329), .O(n2066) );
  NR2P U1995 ( .I1(n1119), .I2(n551), .O(n20) );
  OAI12 U2000 ( .B1(n332), .B2(n2011), .A1(n2012), .O(n896) );
  ND3 U2001 ( .I1(n877), .I2(n2332), .I3(n332), .O(n2012) );
  INV2 U2004 ( .I(n340), .O(n2011) );
  NR2P U2006 ( .I1(n2323), .I2(n499), .O(n2067) );
  BUF2 U2008 ( .I(n1075), .O(n2395) );
  BUF2 U2009 ( .I(n458), .O(n2405) );
  BUF2 U2010 ( .I(n579), .O(n2351) );
  BUF2 U2011 ( .I(n602), .O(n2346) );
  NR2P U2012 ( .I1(decrypt_shift[2]), .I2(decrypt_shift[3]), .O(n1381) );
  BUF2 U2013 ( .I(n515), .O(n2322) );
  OAI12 U2014 ( .B1(n388), .B2(n655), .A1(n2294), .O(n649) );
  ND3 U2015 ( .I1(n655), .I2(n1960), .I3(n388), .O(n2294) );
  ND3 U2016 ( .I1(n768), .I2(n167), .I3(n154), .O(n771) );
  BUF2 U2017 ( .I(n393), .O(n2006) );
  MOAI1 U2018 ( .A1(n13), .A2(n14), .B1(n15), .B2(n16), .O(n11) );
  AO12 U2019 ( .B1(n17), .B2(n18), .A1(n19), .O(n15) );
  BUF2 U2020 ( .I(n393), .O(n2005) );
  OAI112S U2021 ( .C1(n2084), .C2(n2083), .A1(n2085), .B1(n907), .O(n2079) );
  INV2 U2022 ( .I(n1274), .O(n2084) );
  ND3 U2023 ( .I1(n2083), .I2(n2322), .I3(n2086), .O(n2085) );
  NR2 U2024 ( .I1(n916), .I2(n2327), .O(n2086) );
  MOAI1 U2025 ( .A1(n49), .A2(n45), .B1(n44), .B2(n45), .O(n1544) );
  ND3 U2026 ( .I1(n896), .I2(n337), .I3(n323), .O(n2010) );
  NR2 U2027 ( .I1(n2014), .I2(n877), .O(n2013) );
  OAI12S U2028 ( .B1(n332), .B2(n330), .A1(n891), .O(n885) );
  ND3 U2029 ( .I1(n323), .I2(n877), .I3(n892), .O(n891) );
  MOAI1 U2030 ( .A1(n334), .A2(n335), .B1(n336), .B2(n337), .O(n333) );
  OAI12S U2031 ( .B1(n338), .B2(n339), .A1(n330), .O(n336) );
  OAI12S U2032 ( .B1(n2314), .B2(n354), .A1(n363), .O(n360) );
  OAI12S U2033 ( .B1(n1961), .B2(n378), .A1(n383), .O(n391) );
  AOI12S U2034 ( .B1(n319), .B2(n1331), .A1(n342), .O(n1322) );
  ND3 U2035 ( .I1(n378), .I2(n386), .I3(n652), .O(n646) );
  MOAI1 U2036 ( .A1(n653), .A2(n380), .B1(n653), .B2(n654), .O(n652) );
  MOAI1 U2037 ( .A1(n2006), .A2(n1800), .B1(n655), .B2(n656), .O(n654) );
  MOAI1 U2038 ( .A1(n25), .A2(n22), .B1(n21), .B2(n22), .O(n1479) );
  ND3 U2039 ( .I1(n631), .I2(n354), .I3(n366), .O(n625) );
  MOAI1 U2040 ( .A1(n352), .A2(n632), .B1(n632), .B2(n633), .O(n631) );
  MOAI1 U2041 ( .A1(n2314), .A2(n2313), .B1(n634), .B2(n635), .O(n633) );
  MOAI1 U2042 ( .A1(n1917), .A2(n1054), .B1(n1041), .B2(n1044), .O(n1928) );
  BUF1 U2043 ( .I(n220), .O(n2347) );
  BUF1 U2044 ( .I(n829), .O(n2383) );
  ND3 U2045 ( .I1(n388), .I2(n1222), .I3(n648), .O(n1215) );
  AO222 U2046 ( .A1(n1223), .A2(n655), .B1(n1224), .B2(n382), .C1(n650), .C2(
        n653), .O(n1222) );
  NR2 U2047 ( .I1(n653), .I2(n386), .O(n1224) );
  OAI12S U2048 ( .B1(n380), .B2(n645), .A1(n1225), .O(n1223) );
  INV2 U2049 ( .I(encrypt_shift[2]), .O(n2310) );
  AN3B1 U2050 ( .I1(n1332), .I2(n894), .B1(n335), .O(n342) );
  OAI12S U2051 ( .B1(n2292), .B2(n392), .A1(n1800), .O(n2289) );
  AN2 U2052 ( .I1(n378), .I2(n649), .O(n2292) );
  OA22 U2053 ( .A1(n213), .A2(n214), .B1(n215), .B2(n216), .O(n212) );
  AOI13HS U2054 ( .B1(n215), .B2(n217), .B3(n204), .A1(n218), .O(n213) );
  NR2 U2055 ( .I1(n219), .I2(n2348), .O(n218) );
  MAOI1 U2056 ( .A1(n221), .A2(n222), .B1(n223), .B2(n204), .O(n219) );
  OA222 U2057 ( .A1(n382), .A2(n383), .B1(n384), .B2(n385), .C1(n386), .C2(
        n387), .O(n376) );
  ND2 U2058 ( .I1(n1801), .I2(n386), .O(n384) );
  ND2 U2059 ( .I1(n388), .I2(n389), .O(n385) );
  OA12 U2060 ( .B1(n775), .B2(n146), .A1(n165), .O(n770) );
  OA222 U2061 ( .A1(n147), .A2(n776), .B1(n2404), .B2(n777), .C1(n167), .C2(
        n778), .O(n775) );
  ND2 U2062 ( .I1(n779), .I2(n774), .O(n777) );
  XNR2 U2063 ( .I1(n2407), .I2(n2414), .O(n779) );
  AN3B1 U2064 ( .I1(n612), .I2(n613), .B1(n614), .O(n611) );
  INV2 U2065 ( .I(encrypt_shift[4]), .O(n2539) );
  ND2 U2066 ( .I1(n837), .I2(n2383), .O(n830) );
  BUF1 U2067 ( .I(decrypt_shift[4]), .O(n2515) );
  BUF1 U2068 ( .I(decrypt_shift[4]), .O(n2516) );
  BUF1 U2069 ( .I(decrypt_shift[4]), .O(n2513) );
  BUF1 U2070 ( .I(decrypt_shift[4]), .O(n2514) );
  BUF1 U2071 ( .I(n2553), .O(n2543) );
  BUF1 U2072 ( .I(n2553), .O(n2544) );
  BUF1 U2073 ( .I(n2553), .O(n2545) );
  BUF1 U2074 ( .I(n2552), .O(n2548) );
  BUF1 U2075 ( .I(n2552), .O(n2547) );
  BUF1 U2076 ( .I(n2553), .O(n2546) );
  BUF1 U2077 ( .I(n2552), .O(n2549) );
  BUF1 U2078 ( .I(n2552), .O(n2550) );
  BUF1 U2079 ( .I(n2552), .O(n2551) );
  ND2P U2080 ( .I1(decrypt_shift[1]), .I2(decrypt_shift[0]), .O(n2169) );
  ND2P U2081 ( .I1(decrypt_shift[1]), .I2(n2259), .O(n2170) );
  INV2 U2082 ( .I(decrypt_shift[1]), .O(n2260) );
  XNR2P U2083 ( .I1(n1579), .I2(din[18]), .O(n1547) );
  MOAI1 U2084 ( .A1(n2505), .A2(n1580), .B1(n1581), .B2(n2510), .O(n1579) );
  XNR2P U2085 ( .I1(n1582), .I2(din[17]), .O(n49) );
  MOAI1 U2086 ( .A1(n2506), .A2(n1583), .B1(n1584), .B2(n2510), .O(n1582) );
  XOR2P U2087 ( .I1(din[19]), .I2(n1566), .O(n38) );
  MAOI1 U2088 ( .A1(n2498), .A2(n1567), .B1(n2503), .B2(n1568), .O(n1566) );
  XOR2P U2089 ( .I1(din[24]), .I2(n1823), .O(n1002) );
  OA22 U2090 ( .A1(n1824), .A2(n2498), .B1(n2511), .B2(n1825), .O(n1823) );
  XOR2P U2091 ( .I1(din[24]), .I2(n1762), .O(n970) );
  OA22 U2092 ( .A1(n1763), .A2(n2535), .B1(n2529), .B2(n1764), .O(n1762) );
  MOAI1T U2093 ( .A1(n2521), .A2(n2034), .B1(n2035), .B2(n2526), .O(n877) );
  XNR2 U2094 ( .I1(din[24]), .I2(n2036), .O(n2035) );
  XNR2 U2095 ( .I1(n2002), .I2(n1513), .O(n2034) );
  MOAI1T U2096 ( .A1(n2519), .A2(n2122), .B1(n2123), .B2(n2527), .O(n499) );
  XNR2 U2097 ( .I1(din[29]), .I2(n2050), .O(n2123) );
  XNR2 U2098 ( .I1(n2124), .I2(n2040), .O(n2122) );
  MOAI1T U2099 ( .A1(n2527), .A2(n2043), .B1(n2044), .B2(n2526), .O(n337) );
  XNR2 U2100 ( .I1(din[21]), .I2(n1528), .O(n2044) );
  XNR2 U2101 ( .I1(n1994), .I2(n1518), .O(n2043) );
  MOAI1T U2102 ( .A1(n2531), .A2(n2135), .B1(n2136), .B2(n2534), .O(n502) );
  XNR2 U2103 ( .I1(din[27]), .I2(n2130), .O(n2136) );
  XNR2 U2104 ( .I1(n1789), .I2(n1764), .O(n2135) );
  MOAI1T U2105 ( .A1(n2507), .A2(n1660), .B1(n2222), .B2(n2509), .O(n354) );
  XNR2 U2106 ( .I1(din[4]), .I2(n1657), .O(n2222) );
  MOAI1T U2111 ( .A1(n2518), .A2(n1721), .B1(n2300), .B2(n2528), .O(n378) );
  XNR2 U2112 ( .I1(din[4]), .I2(n1718), .O(n2300) );
  MOAI1T U2115 ( .A1(n2517), .A2(n2306), .B1(n2307), .B2(n2523), .O(n386) );
  XNR2 U2117 ( .I1(din[7]), .I2(n1453), .O(n2307) );
  XNR2 U2119 ( .I1(n1898), .I2(n1935), .O(n2306) );
  MOAI1T U2120 ( .A1(n2527), .A2(n1521), .B1(n1522), .B2(n2524), .O(n1119) );
  XNR2 U2121 ( .I1(din[18]), .I2(n1523), .O(n1522) );
  XOR2 U2122 ( .I1(din[18]), .I2(n1524), .O(n1521) );
  MOAI1T U2123 ( .A1(n2521), .A2(n1945), .B1(n1946), .B2(n2526), .O(n613) );
  XNR2 U2124 ( .I1(din[9]), .I2(n1936), .O(n1946) );
  XNR2 U2125 ( .I1(n1893), .I2(n1711), .O(n1945) );
  MOAI1T U2126 ( .A1(n2519), .A2(n2297), .B1(n2298), .B2(n2527), .O(n655) );
  XNR2 U2127 ( .I1(n1881), .I2(n2299), .O(n2297) );
  XNR2 U2128 ( .I1(din[8]), .I2(n1726), .O(n2298) );
  MOAI1T U2129 ( .A1(n2527), .A2(n2046), .B1(n2047), .B2(n2527), .O(n890) );
  XNR2 U2130 ( .I1(n1780), .I2(n1768), .O(n2046) );
  XNR2 U2131 ( .I1(din[23]), .I2(n1515), .O(n2047) );
  MOAI1T U2132 ( .A1(n2531), .A2(n1950), .B1(n1951), .B2(n2534), .O(n1912) );
  XNR2 U2133 ( .I1(din[12]), .I2(n1703), .O(n1951) );
  XNR2 U2134 ( .I1(n1395), .I2(n1722), .O(n1950) );
  MOAI1T U2135 ( .A1(n2522), .A2(n1723), .B1(n1724), .B2(n2524), .O(n837) );
  XNR2 U2136 ( .I1(n1624), .I2(n1726), .O(n1723) );
  XNR2 U2137 ( .I1(din[31]), .I2(n1725), .O(n1724) );
  MOAI1T U2138 ( .A1(n2520), .A2(n1511), .B1(n1512), .B2(n2523), .O(n16) );
  XNR2 U2139 ( .I1(din[19]), .I2(n1513), .O(n1512) );
  XNR2 U2140 ( .I1(n1514), .I2(n1515), .O(n1511) );
  MOAI1T U2141 ( .A1(n2521), .A2(n1525), .B1(n1526), .B2(n2524), .O(n25) );
  XNR2 U2142 ( .I1(din[17]), .I2(n1527), .O(n1526) );
  XOR2 U2143 ( .I1(din[17]), .I2(n1528), .O(n1525) );
  AOI22 U2144 ( .A1(n2504), .A2(n1581), .B1(n1818), .B2(n2512), .O(n1738) );
  MOAI1 U2145 ( .A1(n1372), .A2(n2499), .B1(n1374), .B2(n2503), .O(n1371) );
  AO2222 U2146 ( .A1(n2496), .A2(n1376), .B1(n2493), .B2(n1378), .C1(n2488), 
        .C2(n1380), .D1(n2483), .D2(n1382), .O(n1374) );
  OAI22 U2147 ( .A1(n2511), .A2(n1586), .B1(n1587), .B2(n2504), .O(n1739) );
  MOAI1T U2148 ( .A1(n2521), .A2(n1943), .B1(n1944), .B2(n2526), .O(n1041) );
  XNR2 U2149 ( .I1(n1898), .I2(n1725), .O(n1943) );
  XNR2 U2150 ( .I1(din[7]), .I2(n1701), .O(n1944) );
  MOAI1T U2151 ( .A1(n2520), .A2(n2051), .B1(n2052), .B2(n2527), .O(n894) );
  XNR2 U2152 ( .I1(din[20]), .I2(n2053), .O(n2052) );
  XNR2 U2153 ( .I1(n1519), .I2(n1781), .O(n2051) );
  XOR2 U2154 ( .I1(din[4]), .I2(n2301), .O(n1721) );
  OA2222S U2155 ( .A1(n1952), .A2(n2470), .B1(n1719), .B2(n2474), .C1(n1708), 
        .C2(n1505), .D1(n1707), .D2(n1503), .O(n2301) );
  XNR2 U2156 ( .I1(n1388), .I2(n1468), .O(n1937) );
  XNR2 U2157 ( .I1(din[11]), .I2(n1939), .O(n1938) );
  XOR2 U2158 ( .I1(din[20]), .I2(n1576), .O(n1075) );
  MAOI1 U2159 ( .A1(n1577), .A2(n2506), .B1(n2510), .B2(n1578), .O(n1576) );
  XOR2 U2160 ( .I1(din[25]), .I2(n1773), .O(n723) );
  OA22 U2161 ( .A1(n2529), .A2(n1774), .B1(n1775), .B2(n2532), .O(n1773) );
  OA2222S U2162 ( .A1(n1508), .A2(n2469), .B1(n1506), .B2(n2474), .C1(n1504), 
        .C2(n1505), .D1(n1776), .D2(n1503), .O(n1775) );
  OA2222S U2163 ( .A1(n1776), .A2(n2470), .B1(n1777), .B2(n2474), .C1(n1778), 
        .C2(n1505), .D1(n1510), .D2(n1503), .O(n1774) );
  XOR2 U2164 ( .I1(din[25]), .I2(n1832), .O(n679) );
  OA22 U2165 ( .A1(n2505), .A2(n1833), .B1(n1834), .B2(n2504), .O(n1832) );
  XNR2 U2166 ( .I1(n1899), .I2(din[10]), .O(n579) );
  MOAI1 U2167 ( .A1(n1900), .A2(n2498), .B1(n1901), .B2(n2502), .O(n1899) );
  AO2222 U2168 ( .A1(n2495), .A2(n1380), .B1(n2492), .B2(n1382), .C1(n2487), 
        .C2(n1391), .D1(n2482), .D2(n1392), .O(n1901) );
  XNR2 U2169 ( .I1(n1438), .I2(din[14]), .O(n152) );
  MOAI1 U2170 ( .A1(n1439), .A2(n2530), .B1(n1441), .B2(n2535), .O(n1438) );
  AO2222 U2171 ( .A1(n2479), .A2(n1443), .B1(n2476), .B2(n1445), .C1(n2471), 
        .C2(n1447), .D1(n2466), .D2(n1449), .O(n1441) );
  XNR2 U2172 ( .I1(n1954), .I2(din[10]), .O(n602) );
  MOAI1 U2173 ( .A1(n1955), .A2(n2530), .B1(n1956), .B2(n2534), .O(n1954) );
  AO2222 U2174 ( .A1(n2479), .A2(n1447), .B1(n2476), .B2(n1449), .C1(n2471), 
        .C2(n1457), .D1(n2466), .D2(n1458), .O(n1956) );
  MOAI1P U2175 ( .A1(n2519), .A2(n2131), .B1(n2132), .B2(n2527), .O(n515) );
  XNR2 U2176 ( .I1(din[28]), .I2(n2129), .O(n2132) );
  XNR2 U2177 ( .I1(n1769), .I2(n1530), .O(n2131) );
  MOAI1 U2178 ( .A1(n2548), .A2(n2054), .B1(n2055), .B2(n2552), .O(N1747) );
  XNR2 U2346 ( .I1(din[33]), .I2(n2056), .O(n2055) );
  XOR2 U2347 ( .I1(din[33]), .I2(n2137), .O(n2054) );
  MOAI1T U2348 ( .A1(n2517), .A2(n1450), .B1(n1451), .B2(n2523), .O(n167) );
  XNR2 U2349 ( .I1(din[13]), .I2(n1452), .O(n1451) );
  XNR2 U2350 ( .I1(n1384), .I2(n1453), .O(n1450) );
  XOR2 U2351 ( .I1(din[4]), .I2(n2235), .O(n1660) );
  OA2222S U2352 ( .A1(n1890), .A2(n2486), .B1(n1658), .B2(n2491), .C1(n1647), 
        .C2(n1642), .D1(n1645), .D2(n1640), .O(n2235) );
  MOAI1T U2353 ( .A1(n2531), .A2(n2127), .B1(n2128), .B2(n2534), .O(n916) );
  XNR2 U2354 ( .I1(n1624), .I2(n2130), .O(n2127) );
  XNR2 U2355 ( .I1(din[31]), .I2(n2129), .O(n2128) );
  MOAI1P U2356 ( .A1(n2520), .A2(n2048), .B1(n2049), .B2(n2525), .O(n1320) );
  XNR2 U2357 ( .I1(n1997), .I2(n2050), .O(n2048) );
  XNR2 U2358 ( .I1(din[22]), .I2(n1790), .O(n2049) );
  MOAI1P U2359 ( .A1(n2520), .A2(n1755), .B1(n1756), .B2(n2525), .O(n708) );
  XOR2 U2360 ( .I1(din[26]), .I2(n1523), .O(n1755) );
  XNR2 U2361 ( .I1(din[26]), .I2(n1757), .O(n1756) );
  MOAI1P U2362 ( .A1(n2521), .A2(n1695), .B1(n1696), .B2(n2524), .O(n280) );
  XNR2 U2363 ( .I1(din[1]), .I2(n1469), .O(n1696) );
  XNR2 U2364 ( .I1(n1630), .I2(n1701), .O(n1695) );
  MOAI1P U2365 ( .A1(n2518), .A2(n1466), .B1(n1467), .B2(n2523), .O(n458) );
  XNR2 U2366 ( .I1(din[15]), .I2(n1468), .O(n1467) );
  XNR2 U2367 ( .I1(n1402), .I2(n1469), .O(n1466) );
  MOAI1P U2368 ( .A1(n2522), .A2(n1933), .B1(n1934), .B2(n2525), .O(n220) );
  XNR2 U2369 ( .I1(n1881), .I2(n1936), .O(n1933) );
  XNR2 U2370 ( .I1(din[8]), .I2(n1935), .O(n1934) );
  MOAI1P U2371 ( .A1(n2520), .A2(n1516), .B1(n1517), .B2(n2524), .O(n1104) );
  XNR2 U2372 ( .I1(din[20]), .I2(n1518), .O(n1517) );
  XNR2 U2373 ( .I1(n1519), .I2(n1520), .O(n1516) );
  MOAI1P U2374 ( .A1(n2522), .A2(n1709), .B1(n1710), .B2(n2524), .O(n829) );
  XNR2 U2375 ( .I1(din[0]), .I2(n1711), .O(n1710) );
  XNR2 U2376 ( .I1(n1649), .I2(n1464), .O(n1709) );
  MOAI1P U2377 ( .A1(n2526), .A2(n2038), .B1(n2039), .B2(n2525), .O(n889) );
  XNR2 U2378 ( .I1(n1514), .I2(n1527), .O(n2038) );
  XNR2 U2379 ( .I1(din[19]), .I2(n2040), .O(n2039) );
  MOAI1P U2380 ( .A1(n2518), .A2(n2302), .B1(n2303), .B2(n2528), .O(n393) );
  XNR2 U2381 ( .I1(din[6]), .I2(n1455), .O(n2303) );
  XNR2 U2382 ( .I1(n2253), .I2(n1955), .O(n2302) );
  MOAI1P U2383 ( .A1(n2518), .A2(n1462), .B1(n1463), .B2(n2523), .O(n144) );
  XNR2 U2384 ( .I1(n1398), .I2(n1465), .O(n1462) );
  XNR2 U2385 ( .I1(din[16]), .I2(n1464), .O(n1463) );
  MOAI1P U2386 ( .A1(n2522), .A2(n1783), .B1(n1784), .B2(n2526), .O(n59) );
  XNR2 U2387 ( .I1(din[27]), .I2(n1520), .O(n1784) );
  XNR2 U2388 ( .I1(n1789), .I2(n1790), .O(n1783) );
  MOAI1P U2389 ( .A1(n2523), .A2(n1766), .B1(n1767), .B2(n2525), .O(n66) );
  XNR2 U2390 ( .I1(din[28]), .I2(n1768), .O(n1767) );
  XNR2 U2391 ( .I1(n1769), .I2(n1757), .O(n1766) );
  MOAI1P U2392 ( .A1(n2517), .A2(n2308), .B1(n2309), .B2(n2525), .O(n390) );
  XNR2 U2393 ( .I1(n1637), .I2(n1452), .O(n2308) );
  XNR2 U2394 ( .I1(din[3]), .I2(n1465), .O(n2309) );
  MOAI1P U2395 ( .A1(n2517), .A2(n2304), .B1(n2305), .B2(n2527), .O(n377) );
  XNR2 U2396 ( .I1(din[5]), .I2(n2299), .O(n2305) );
  XNR2 U2397 ( .I1(n2255), .I2(n1939), .O(n2304) );
  MOAI1P U2398 ( .A1(n2519), .A2(n2125), .B1(n2126), .B2(n2528), .O(n496) );
  XNR2 U2399 ( .I1(n1649), .I2(n2053), .O(n2125) );
  XNR2 U2400 ( .I1(din[0]), .I2(n1501), .O(n2126) );
  XOR2 U2401 ( .I1(din[2]), .I2(n1655), .O(n813) );
  OA22 U2402 ( .A1(n1656), .A2(n2498), .B1(n2512), .B2(n1657), .O(n1655) );
  OA2222S U2403 ( .A1(n1658), .A2(n2486), .B1(n1647), .B2(n2491), .C1(n1645), 
        .C2(n1642), .D1(n1643), .D2(n1640), .O(n1656) );
  XOR2 U2404 ( .I1(din[2]), .I2(n1716), .O(n836) );
  OA22 U2405 ( .A1(n1717), .A2(n2535), .B1(n2529), .B2(n1718), .O(n1716) );
  OA2222S U2406 ( .A1(n1719), .A2(n2470), .B1(n1708), .B2(n2474), .C1(n1707), 
        .C2(n1505), .D1(n1706), .D2(n1503), .O(n1717) );
  XOR2 U2407 ( .I1(din[27]), .I2(n1841), .O(n85) );
  OA22 U2408 ( .A1(n2511), .A2(n1842), .B1(n1578), .B2(n2499), .O(n1841) );
  MOAI1P U2409 ( .A1(n2520), .A2(n2087), .B1(n2088), .B2(n2528), .O(n514) );
  XNR2 U2410 ( .I1(din[30]), .I2(n1524), .O(n2088) );
  XNR2 U2411 ( .I1(n2105), .I2(n2036), .O(n2087) );
  INV2 U2412 ( .I(din[24]), .O(n2002) );
  INV2 U2413 ( .I(din[31]), .O(n1624) );
  INV2 U2414 ( .I(din[28]), .O(n1769) );
  INV2 U2415 ( .I(din[8]), .O(n1881) );
  INV2 U2416 ( .I(din[7]), .O(n1898) );
  INV2 U2417 ( .I(din[12]), .O(n1395) );
  INV2 U2418 ( .I(din[23]), .O(n1780) );
  INV2 U2419 ( .I(din[0]), .O(n1649) );
  INV2 U2420 ( .I(din[15]), .O(n1402) );
  INV2 U2421 ( .I(din[3]), .O(n1637) );
  INV2 U2422 ( .I(din[19]), .O(n1514) );
  INV2 U2423 ( .I(din[16]), .O(n1398) );
  INV2 U2424 ( .I(din[27]), .O(n1789) );
  INV2 U2425 ( .I(din[20]), .O(n1519) );
  INV2 U2426 ( .I(din[4]), .O(n1661) );
  INV2 U2427 ( .I(din[22]), .O(n1997) );
  INV2 U2428 ( .I(din[6]), .O(n2253) );
  INV2 U2429 ( .I(din[9]), .O(n1893) );
  INV2 U2430 ( .I(din[13]), .O(n1384) );
  INV2 U2431 ( .I(din[1]), .O(n1630) );
  INV2 U2432 ( .I(din[5]), .O(n2255) );
  INV2 U2433 ( .I(din[30]), .O(n2105) );
  INV2 U2434 ( .I(din[29]), .O(n2124) );
  INV2 U2435 ( .I(din[21]), .O(n1994) );
  BUF1 U2436 ( .I(n2554), .O(n2553) );
  INV2 U2437 ( .I(stall), .O(N1778) );
  MOAI1 U2438 ( .A1(n2541), .A2(n287), .B1(n288), .B2(n2542), .O(N1772) );
  XOR2 U2439 ( .I1(din[58]), .I2(n316), .O(n287) );
  XNR2 U2440 ( .I1(din[58]), .I2(n289), .O(n288) );
  MOAI1 U2441 ( .A1(n2541), .A2(n843), .B1(n844), .B2(n2540), .O(N1762) );
  XNR2 U2442 ( .I1(din[48]), .I2(n872), .O(n843) );
  XOR2 U2443 ( .I1(n845), .I2(din[48]), .O(n844) );
  MOAI1 U2444 ( .A1(n2540), .A2(n2182), .B1(n2183), .B2(n2542), .O(N1746) );
  XNR2 U2445 ( .I1(din[32]), .I2(n2261), .O(n2182) );
  XOR2 U2446 ( .I1(n2184), .I2(din[32]), .O(n2183) );
  MOAI1 U2447 ( .A1(n2548), .A2(n1727), .B1(n1728), .B2(n2550), .O(N1750) );
  XNR2 U2448 ( .I1(din[36]), .I2(n1729), .O(n1728) );
  XOR2 U2449 ( .I1(din[36]), .I2(n1791), .O(n1727) );
  MOAI1 U2450 ( .A1(n2547), .A2(n1470), .B1(n1471), .B2(n2549), .O(N1752) );
  XOR2 U2451 ( .I1(n1472), .I2(din[38]), .O(n1471) );
  XNR2 U2452 ( .I1(din[38]), .I2(n1536), .O(n1470) );
  MOAI1 U2453 ( .A1(n2546), .A2(n940), .B1(n941), .B2(n2549), .O(N1760) );
  XOR2 U2454 ( .I1(n942), .I2(din[46]), .O(n941) );
  XNR2 U2455 ( .I1(din[46]), .I2(n974), .O(n940) );
  MOAI1 U2456 ( .A1(n2546), .A2(n899), .B1(n900), .B2(n2550), .O(N1761) );
  XOR2 U2457 ( .I1(n901), .I2(din[47]), .O(n900) );
  XNR2 U2458 ( .I1(din[47]), .I2(n921), .O(n899) );
  MOAI1 U2459 ( .A1(n2545), .A2(n52), .B1(n53), .B2(n2551), .O(N1776) );
  XOR2 U2460 ( .I1(n54), .I2(din[62]), .O(n53) );
  XNR2 U2461 ( .I1(din[62]), .I2(n81), .O(n52) );
  MOAI1 U2462 ( .A1(n2547), .A2(n3), .B1(n4), .B2(n2551), .O(N1777) );
  XNR2 U2463 ( .I1(din[63]), .I2(n28), .O(n3) );
  XOR2 U2464 ( .I1(n5), .I2(din[63]), .O(n4) );
  MOAI1 U2465 ( .A1(n2541), .A2(n795), .B1(n796), .B2(n2542), .O(N1763) );
  XNR2 U2466 ( .I1(din[49]), .I2(n820), .O(n795) );
  XOR2 U2467 ( .I1(n797), .I2(din[49]), .O(n796) );
  MOAI1 U2468 ( .A1(n2541), .A2(n519), .B1(n520), .B2(n2542), .O(N1768) );
  XNR2 U2469 ( .I1(din[54]), .I2(n544), .O(n519) );
  XOR2 U2470 ( .I1(n521), .I2(din[54]), .O(n520) );
  MOAI1 U2471 ( .A1(n2541), .A2(n397), .B1(n398), .B2(n2542), .O(N1770) );
  XNR2 U2472 ( .I1(din[56]), .I2(n431), .O(n397) );
  XOR2 U2473 ( .I1(n399), .I2(din[56]), .O(n398) );
  MOAI1 U2474 ( .A1(n2540), .A2(n1957), .B1(n1958), .B2(encrypt_in), .O(N1748)
         );
  XNR2 U2475 ( .I1(din[34]), .I2(n2004), .O(n1957) );
  XOR2 U2476 ( .I1(n1959), .I2(din[34]), .O(n1958) );
  MOAI1 U2477 ( .A1(n2540), .A2(n1847), .B1(n1848), .B2(n2540), .O(N1749) );
  XOR2 U2478 ( .I1(din[35]), .I2(n1902), .O(n1847) );
  XNR2 U2479 ( .I1(din[35]), .I2(n1849), .O(n1848) );
  MOAI1 U2480 ( .A1(n2540), .A2(n1333), .B1(n1334), .B2(n2540), .O(N1753) );
  XOR2 U2481 ( .I1(din[39]), .I2(n1405), .O(n1333) );
  XNR2 U2482 ( .I1(din[39]), .I2(n1335), .O(n1334) );
  MOAI1 U2483 ( .A1(n2540), .A2(n1279), .B1(n1280), .B2(n2540), .O(N1754) );
  XOR2 U2484 ( .I1(din[40]), .I2(n1308), .O(n1279) );
  XNR2 U2485 ( .I1(din[40]), .I2(n1281), .O(n1280) );
  MOAI1 U2486 ( .A1(n2541), .A2(n1226), .B1(n1227), .B2(n2540), .O(N1755) );
  XOR2 U2487 ( .I1(din[41]), .I2(n1253), .O(n1226) );
  XNR2 U2488 ( .I1(din[41]), .I2(n1228), .O(n1227) );
  MOAI1 U2489 ( .A1(n2541), .A2(n1177), .B1(n1178), .B2(n2542), .O(N1756) );
  XOR2 U2490 ( .I1(din[42]), .I2(n1202), .O(n1177) );
  XNR2 U2491 ( .I1(din[42]), .I2(n1179), .O(n1178) );
  MOAI1 U2492 ( .A1(n2541), .A2(n1121), .B1(n1122), .B2(n2542), .O(N1757) );
  XOR2 U2493 ( .I1(din[43]), .I2(n1150), .O(n1121) );
  XNR2 U2494 ( .I1(din[43]), .I2(n1123), .O(n1122) );
  MOAI1 U2495 ( .A1(n2541), .A2(n1006), .B1(n1007), .B2(n2540), .O(N1759) );
  XOR2 U2496 ( .I1(din[45]), .I2(n1033), .O(n1006) );
  XNR2 U2497 ( .I1(din[45]), .I2(n1008), .O(n1007) );
  MOAI1 U2498 ( .A1(n2541), .A2(n616), .B1(n617), .B2(n2542), .O(N1766) );
  XOR2 U2499 ( .I1(din[52]), .I2(n639), .O(n616) );
  XNR2 U2500 ( .I1(din[52]), .I2(n618), .O(n617) );
  MOAI1 U2501 ( .A1(n2541), .A2(n568), .B1(n569), .B2(n2542), .O(N1767) );
  XOR2 U2502 ( .I1(din[53]), .I2(n593), .O(n568) );
  XNR2 U2503 ( .I1(din[53]), .I2(n570), .O(n569) );
  MOAI1 U2504 ( .A1(n2541), .A2(n343), .B1(n344), .B2(n2542), .O(N1771) );
  XNR2 U2505 ( .I1(din[57]), .I2(n371), .O(n343) );
  XNR2 U2506 ( .I1(din[57]), .I2(n345), .O(n344) );
  MOAI1 U2507 ( .A1(n2540), .A2(n229), .B1(n230), .B2(n2542), .O(N1773) );
  XOR2 U2508 ( .I1(din[59]), .I2(n259), .O(n229) );
  XNR2 U2509 ( .I1(din[59]), .I2(n231), .O(n230) );
  MOAI1 U2510 ( .A1(n2540), .A2(n171), .B1(n172), .B2(n2542), .O(N1774) );
  XOR2 U2511 ( .I1(din[60]), .I2(n201), .O(n171) );
  XNR2 U2512 ( .I1(din[60]), .I2(n173), .O(n172) );
  MOAI1 U2513 ( .A1(n2540), .A2(n108), .B1(n109), .B2(encrypt_in), .O(N1775)
         );
  XNR2 U2514 ( .I1(din[61]), .I2(n140), .O(n108) );
  XNR2 U2515 ( .I1(din[61]), .I2(n110), .O(n109) );
  MOAI1 U2516 ( .A1(n2541), .A2(n462), .B1(n463), .B2(n2542), .O(N1769) );
  XNR2 U2517 ( .I1(din[55]), .I2(n492), .O(n462) );
  XOR2 U2518 ( .I1(n464), .I2(din[55]), .O(n463) );
  INV2 U2519 ( .I(key_in[37]), .O(n2115) );
  INV2 U2520 ( .I(key_in[4]), .O(n2119) );
  INV2 U2521 ( .I(key_in[7]), .O(n2091) );
  INV2 U2522 ( .I(key_in[6]), .O(n2102) );
  INV2 U2523 ( .I(key_in[38]), .O(n2107) );
  INV2 U2524 ( .I(key_in[29]), .O(n2116) );
  INV2 U2525 ( .I(key_in[61]), .O(n2120) );
  INV2 U2526 ( .I(key_in[31]), .O(n2099) );
  INV2 U2527 ( .I(key_in[30]), .O(n2108) );
  INV2 U2528 ( .I(key_in[45]), .O(n2114) );
  INV2 U2529 ( .I(key_in[47]), .O(n2097) );
  INV2 U2530 ( .I(key_in[15]), .O(n2089) );
  INV2 U2531 ( .I(key_in[12]), .O(n2118) );
  INV2 U2532 ( .I(key_in[46]), .O(n2106) );
  INV2 U2533 ( .I(key_in[5]), .O(n2111) );
  INV2 U2534 ( .I(key_in[62]), .O(n2112) );
  INV2 U2535 ( .I(key_in[21]), .O(n2117) );
  INV2 U2536 ( .I(key_in[20]), .O(n2095) );
  INV2 U2537 ( .I(key_in[54]), .O(n2113) );
  MOAI1 U2538 ( .A1(n2541), .A2(n1058), .B1(n1059), .B2(n2542), .O(N1758) );
  XNR2 U2539 ( .I1(din[44]), .I2(n1089), .O(n1058) );
  XOR2 U2540 ( .I1(n1060), .I2(din[44]), .O(n1059) );
  MOAI1 U2541 ( .A1(n2540), .A2(n1592), .B1(n1593), .B2(n2540), .O(N1751) );
  XNR2 U2542 ( .I1(din[37]), .I2(n1663), .O(n1592) );
  XOR2 U2543 ( .I1(n1594), .I2(din[37]), .O(n1593) );
  INV2 U2544 ( .I(key_in[13]), .O(n2110) );
  INV2 U2545 ( .I(key_in[53]), .O(n2121) );
  INV2 U2546 ( .I(key_in[55]), .O(n2104) );
  INV2 U2547 ( .I(key_in[63]), .O(n2103) );
  INV2 U2548 ( .I(key_in[28]), .O(n2093) );
  INV2 U2549 ( .I(key_in[22]), .O(n2109) );
  MOAI1 U2550 ( .A1(n2541), .A2(n730), .B1(n731), .B2(n2542), .O(N1764) );
  XOR2 U2551 ( .I1(din[50]), .I2(n764), .O(n730) );
  XNR2 U2552 ( .I1(din[50]), .I2(n732), .O(n731) );
  MOAI1 U2553 ( .A1(n2541), .A2(n660), .B1(n661), .B2(n2542), .O(N1765) );
  XOR2 U2554 ( .I1(din[51]), .I2(n696), .O(n660) );
  XNR2 U2555 ( .I1(din[51]), .I2(n662), .O(n661) );
  INV2 U2556 ( .I(key_in[44]), .O(n2230) );
  INV2 U2557 ( .I(key_in[42]), .O(n2243) );
  INV2 U2558 ( .I(key_in[41]), .O(n2251) );
  INV2 U2559 ( .I(key_in[25]), .O(n2232) );
  INV2 U2560 ( .I(key_in[59]), .O(n2224) );
  INV2 U2561 ( .I(key_in[60]), .O(n2228) );
  INV2 U2562 ( .I(key_in[57]), .O(n2249) );
  INV2 U2563 ( .I(key_in[58]), .O(n2241) );
  INV2 U2564 ( .I(key_in[26]), .O(n2245) );
  INV2 U2565 ( .I(key_in[27]), .O(n2237) );
  INV2 U2566 ( .I(key_in[17]), .O(n2233) );
  INV2 U2567 ( .I(key_in[50]), .O(n2242) );
  INV2 U2568 ( .I(key_in[18]), .O(n2246) );
  INV2 U2569 ( .I(key_in[36]), .O(n2223) );
  INV2 U2570 ( .I(key_in[1]), .O(n2227) );
  INV2 U2571 ( .I(key_in[2]), .O(n2248) );
  INV2 U2572 ( .I(key_in[39]), .O(n2098) );
  INV2 U2573 ( .I(key_in[14]), .O(n2101) );
  INV2 U2574 ( .I(key_in[23]), .O(n2100) );
  INV2 U2575 ( .I(key_in[33]), .O(n2231) );
  INV2 U2576 ( .I(key_in[51]), .O(n2225) );
  INV2 U2577 ( .I(key_in[52]), .O(n2229) );
  INV2 U2578 ( .I(key_in[9]), .O(n2234) );
  INV2 U2579 ( .I(key_in[43]), .O(n2226) );
  INV2 U2580 ( .I(key_in[49]), .O(n2250) );
  INV2 U2581 ( .I(key_in[3]), .O(n2240) );
  INV2 U2582 ( .I(key_in[34]), .O(n2244) );
  INV2 U2583 ( .I(key_in[10]), .O(n2247) );
  INV2 U2584 ( .I(key_in[35]), .O(n2236) );
  INV2 U2585 ( .I(key_in[19]), .O(n2238) );
  INV2 U2586 ( .I(key_in[11]), .O(n2239) );
  INV2 U2587 ( .I(encrypt_in), .O(n2554) );
  BUF1 U2588 ( .I(test_mode), .O(n2555) );
  XOR2T U2589 ( .I1(n1648), .I2(n1649), .O(n806) );
  QDFZRBS dout_reg_62 ( .D(din[30]), .TD(dout[61]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[62]) );
  QDFZRBS dout_reg_61 ( .D(din[29]), .TD(dout[60]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[61]) );
  QDFZRBS dout_reg_58 ( .D(din[26]), .TD(dout[57]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[58]) );
  QDFZRBS dout_reg_57 ( .D(din[25]), .TD(dout[56]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[57]) );
  QDFZRBS dout_reg_53 ( .D(din[21]), .TD(dout[52]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[53]) );
  QDFZRBS dout_reg_51 ( .D(din[19]), .TD(dout[50]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[51]) );
  QDFZRBS dout_reg_50 ( .D(din[18]), .TD(dout[49]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[50]) );
  QDFZRBS dout_reg_49 ( .D(din[17]), .TD(dout[48]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[49]) );
  QDFZRBS dout_reg_47 ( .D(din[15]), .TD(dout[46]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[47]) );
  QDFZRBS dout_reg_46 ( .D(din[14]), .TD(dout[45]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[46]) );
  QDFZRBS dout_reg_42 ( .D(din[10]), .TD(dout[41]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[42]) );
  QDFZRBS dout_reg_41 ( .D(din[9]), .TD(dout[40]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[41]) );
  QDFZRBS dout_reg_38 ( .D(din[6]), .TD(dout[37]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[38]) );
  QDFZRBS dout_reg_37 ( .D(din[5]), .TD(dout[36]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[37]) );
  QDFZRBS dout_reg_35 ( .D(din[3]), .TD(dout[34]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[35]) );
  QDFZRBS dout_reg_34 ( .D(din[2]), .TD(dout[33]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[34]) );
  QDFZRBS dout_reg_33 ( .D(din[1]), .TD(dout[32]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[33]) );
  QDFZRBS dout_reg_31 ( .D(N1777), .TD(dout[30]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[31]) );
  QDFZRBS dout_reg_30 ( .D(N1776), .TD(dout[29]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[30]) );
  QDFZRBS dout_reg_29 ( .D(N1775), .TD(dout[28]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[29]) );
  QDFZRBS dout_reg_28 ( .D(N1774), .TD(dout[27]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[28]) );
  QDFZRBS dout_reg_27 ( .D(N1773), .TD(dout[26]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[27]) );
  QDFZRBS dout_reg_26 ( .D(N1772), .TD(dout[25]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[26]) );
  QDFZRBS dout_reg_25 ( .D(N1771), .TD(dout[24]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[25]) );
  QDFZRBS dout_reg_23 ( .D(N1769), .TD(dout[22]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[23]) );
  QDFZRBS dout_reg_21 ( .D(N1767), .TD(dout[20]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[21]) );
  QDFZRBS dout_reg_20 ( .D(N1766), .TD(dout[19]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[20]) );
  QDFZRBS dout_reg_19 ( .D(N1765), .TD(dout[18]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[19]) );
  QDFZRBS dout_reg_18 ( .D(N1764), .TD(dout[17]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[18]) );
  QDFZRBS dout_reg_17 ( .D(N1763), .TD(dout[16]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[17]) );
  QDFZRBS dout_reg_16 ( .D(N1762), .TD(dout[15]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[16]) );
  QDFZRBS dout_reg_15 ( .D(N1761), .TD(dout[14]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[15]) );
  QDFZRBS dout_reg_14 ( .D(N1760), .TD(dout[13]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[14]) );
  QDFZRBS dout_reg_13 ( .D(N1759), .TD(dout[12]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[13]) );
  QDFZRBS dout_reg_12 ( .D(N1758), .TD(dout[11]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[12]) );
  QDFZRBS dout_reg_11 ( .D(N1757), .TD(dout[10]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[11]) );
  QDFZRBS dout_reg_10 ( .D(N1756), .TD(dout[9]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[10]) );
  QDFZRBS dout_reg_8 ( .D(N1754), .TD(dout[7]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[8]) );
  QDFZRBS dout_reg_7 ( .D(N1753), .TD(dout[6]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[7]) );
  QDFZRBS dout_reg_6 ( .D(N1752), .TD(dout[5]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[6]) );
  QDFZRBS dout_reg_5 ( .D(N1751), .TD(dout[4]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[5]) );
  QDFZRBS dout_reg_4 ( .D(N1750), .TD(dout[3]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[4]) );
  QDFZRBS dout_reg_3 ( .D(N1749), .TD(dout[2]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[3]) );
  QDFZRBS dout_reg_2 ( .D(N1748), .TD(dout[1]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[2]) );
  QDFZRBS dout_reg_1 ( .D(N1747), .TD(dout[0]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[1]) );
  QDFZRBS dout_reg_0 ( .D(N1746), .TD(n2557), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[0]) );
  QDFZRBS dout_reg_9 ( .D(N1755), .TD(dout[8]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[9]) );
  QDFZRBS dout_reg_63 ( .D(din[31]), .TD(dout[62]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[63]) );
  QDFZRBS dout_reg_60 ( .D(din[28]), .TD(dout[59]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[60]) );
  QDFZRBS dout_reg_59 ( .D(din[27]), .TD(dout[58]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[59]) );
  QDFZRBS dout_reg_56 ( .D(din[24]), .TD(dout[55]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[56]) );
  QDFZRBS dout_reg_55 ( .D(din[23]), .TD(dout[54]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[55]) );
  QDFZRBS dout_reg_54 ( .D(din[22]), .TD(dout[53]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[54]) );
  QDFZRBS dout_reg_52 ( .D(din[20]), .TD(dout[51]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[52]) );
  QDFZRBS dout_reg_48 ( .D(din[16]), .TD(dout[47]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[48]) );
  QDFZRBS dout_reg_45 ( .D(din[13]), .TD(dout[44]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[45]) );
  QDFZRBS dout_reg_44 ( .D(din[12]), .TD(dout[43]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[44]) );
  QDFZRBS dout_reg_43 ( .D(din[11]), .TD(dout[42]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[43]) );
  QDFZRBS dout_reg_40 ( .D(din[8]), .TD(dout[39]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[40]) );
  QDFZRBS dout_reg_39 ( .D(din[7]), .TD(dout[38]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[39]) );
  QDFZRBS dout_reg_36 ( .D(din[4]), .TD(dout[35]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[36]) );
  QDFZRBS dout_reg_32 ( .D(din[0]), .TD(dout[31]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[32]) );
  QDFZRBS dout_reg_24 ( .D(N1770), .TD(dout[23]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[24]) );
  QDFZRBS dout_reg_22 ( .D(N1768), .TD(dout[21]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N1778_0_0), .RB(POR), .Q(dout[22]) );
endmodule


module tiny_des ( hclk, POR, hresetn, encrypt, edr, key_in, din, din_valid, 
        round, dout, dout_valid, test_mode, test_se, test_si );
  input [1:0] edr;
  input [63:0] key_in;
  input [63:0] din;
  output [3:0] round;
  output [63:0] dout;
  input hclk, POR, hresetn, encrypt, din_valid, test_mode, test_se, test_si;
  output dout_valid;
  wire   n87, state, N37, N38, N39, N40, stall, N66, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n1, n2, n4, n5, n6, n7, n8,
         n9, n10, n61, n81, n82, n83, n84, n85, n86;
  wire   [63:0] r_din;
  wire   [4:0] encrypt_shift;
  wire   [4:0] decrypt_shift;

  AO22P U23 ( .A1(dout[24]), .A2(n7), .B1(din[25]), .B2(n83), .O(r_din[4]) );
  AO22P U51 ( .A1(dout[62]), .A2(n5), .B1(din[63]), .B2(n10), .O(r_din[24]) );
  OR3B2P U82 ( .I1(encrypt_shift[4]), .B1(n37), .B2(n38), .O(encrypt_shift[0])
         );
  tiny_des_round u_tiny_des_round ( .hclk(hclk), .POR(POR), .hresetn(hresetn), 
        .stall(stall), .encrypt_in(encrypt), .encrypt_shift(encrypt_shift), 
        .decrypt_shift(decrypt_shift), .key_in(key_in), .din(r_din), .dout({
        dout[7], dout[15], dout[23], dout[31], dout[39], dout[47], dout[55], 
        dout[63], dout[5], dout[13], dout[21], dout[29], dout[37], dout[45], 
        dout[53], dout[61], dout[3], dout[11], dout[19], dout[27], dout[35], 
        dout[43], dout[51], dout[59], dout[1], dout[9], dout[17], dout[25], 
        dout[33], dout[41], dout[49], dout[57], dout[6], dout[14], dout[22], 
        dout[30], dout[38], dout[46], dout[54], dout[62], dout[4], dout[12], 
        dout[20], dout[28], dout[36], dout[44], dout[52], dout[60], dout[2], 
        dout[10], dout[18], dout[26], dout[34], dout[42], dout[50], dout[58], 
        dout[0], dout[8], dout[16], dout[24], dout[32], dout[40], dout[48], 
        dout[56]}), .test_mode(test_mode), .test_se(test_se), .test_si(state)
         );
  AO22 U3 ( .A1(dout[56]), .A2(n4), .B1(din[57]), .B2(n8), .O(r_din[0]) );
  AO22 U4 ( .A1(dout[0]), .A2(n4), .B1(din[1]), .B2(n85), .O(r_din[7]) );
  AO22 U5 ( .A1(dout[58]), .A2(n4), .B1(din[59]), .B2(n85), .O(r_din[8]) );
  AO22 U6 ( .A1(dout[60]), .A2(n4), .B1(din[61]), .B2(n9), .O(r_din[16]) );
  AO22 U7 ( .A1(dout[28]), .A2(n5), .B1(din[29]), .B2(n10), .O(r_din[20]) );
  AO22 U8 ( .A1(dout[38]), .A2(n5), .B1(din[39]), .B2(n61), .O(r_din[27]) );
  AO22 U9 ( .A1(dout[30]), .A2(n5), .B1(din[31]), .B2(n61), .O(r_din[28]) );
  AO22 U10 ( .A1(dout[6]), .A2(n5), .B1(din[7]), .B2(n61), .O(r_din[31]) );
  AO22 U11 ( .A1(dout[52]), .A2(n4), .B1(din[53]), .B2(n9), .O(r_din[17]) );
  AO22 U12 ( .A1(dout[44]), .A2(n5), .B1(din[45]), .B2(n9), .O(r_din[18]) );
  AO22 U13 ( .A1(dout[36]), .A2(n4), .B1(din[37]), .B2(n9), .O(r_din[19]) );
  AO22 U14 ( .A1(dout[46]), .A2(n5), .B1(din[47]), .B2(n10), .O(r_din[26]) );
  ND3 U15 ( .I1(round[2]), .I2(round[3]), .I3(n58), .O(n40) );
  ND3P U16 ( .I1(round[2]), .I2(round[3]), .I3(n56), .O(n24) );
  ND3P U17 ( .I1(round[2]), .I2(round[3]), .I3(n50), .O(n25) );
  INV1 U18 ( .I(n28), .O(n46) );
  ND3 U19 ( .I1(n49), .I2(n55), .I3(n34), .O(n27) );
  OAI112 U20 ( .C1(n20), .C2(n29), .A1(n30), .B1(n31), .O(encrypt_shift[2]) );
  ND2 U21 ( .I1(round[0]), .I2(n23), .O(n47) );
  OAI112 U22 ( .C1(n47), .C2(n20), .A1(n30), .B1(n48), .O(decrypt_shift[2]) );
  OR3B2 U24 ( .I1(n1), .B1(n43), .B2(n62), .O(decrypt_shift[0]) );
  OAI22 U25 ( .A1(n69), .A2(n36), .B1(n18), .B2(n29), .O(n1) );
  ND3P U26 ( .I1(n24), .I2(n25), .I3(n26), .O(encrypt_shift[3]) );
  ND3P U27 ( .I1(n46), .I2(n20), .I3(n45), .O(decrypt_shift[3]) );
  NR2P U28 ( .I1(round[1]), .I2(round[0]), .O(n58) );
  NR2P U29 ( .I1(n18), .I2(round[3]), .O(n68) );
  ND2P U30 ( .I1(round[3]), .I2(n18), .O(n20) );
  INV2 U31 ( .I(n27), .O(n43) );
  INV3 U32 ( .I(n8), .O(n4) );
  ND2 U33 ( .I1(n37), .I2(n57), .O(n28) );
  NR2P U34 ( .I1(n65), .I2(n53), .O(n33) );
  INV2 U35 ( .I(n47), .O(n50) );
  ND2P U36 ( .I1(n35), .I2(n36), .O(encrypt_shift[1]) );
  NR2P U37 ( .I1(n50), .I2(n56), .O(n42) );
  INV2 U38 ( .I(n38), .O(n59) );
  INV2 U39 ( .I(n56), .O(n53) );
  INV3 U40 ( .I(n8), .O(n5) );
  NR2 U41 ( .I1(n42), .I2(n75), .O(N38) );
  BUF2 U42 ( .I(n86), .O(n8) );
  OA112 U43 ( .C1(n53), .C2(n20), .A1(n30), .B1(n54), .O(n35) );
  AN2 U44 ( .I1(n24), .I2(n55), .O(n54) );
  AN3 U45 ( .I1(n40), .I2(n44), .I3(n46), .O(n30) );
  OR2B1 U46 ( .I1(n20), .B1(n58), .O(n37) );
  OA112 U47 ( .C1(n38), .C2(n21), .A1(n25), .B1(n49), .O(n48) );
  NR2T U48 ( .I1(n23), .I2(round[0]), .O(n56) );
  AOI112P U49 ( .C1(n63), .C2(n59), .A1(n64), .B1(n33), .O(n62) );
  INV2 U50 ( .I(n44), .O(n64) );
  ND2P U52 ( .I1(n66), .I2(n50), .O(n36) );
  ND2P U53 ( .I1(n66), .I2(n58), .O(n38) );
  ND3 U54 ( .I1(n39), .I2(n40), .I3(n41), .O(encrypt_shift[4]) );
  AO12 U55 ( .B1(n29), .B2(n42), .A1(n20), .O(n39) );
  AN2 U56 ( .I1(n25), .I2(n24), .O(n41) );
  ND2P U57 ( .I1(n66), .I2(n67), .O(n44) );
  ND2 U58 ( .I1(n67), .I2(n68), .O(n57) );
  ND2 U59 ( .I1(n68), .I2(n56), .O(n34) );
  INV2 U60 ( .I(n29), .O(n67) );
  ND2 U61 ( .I1(n68), .I2(n58), .O(n49) );
  ND2 U62 ( .I1(n68), .I2(n50), .O(n55) );
  INV2 U63 ( .I(n66), .O(n65) );
  NR2 U64 ( .I1(n32), .I2(n33), .O(n31) );
  INV2 U65 ( .I(n34), .O(n32) );
  INV2 U66 ( .I(n13), .O(n63) );
  NR2 U67 ( .I1(n27), .I2(n28), .O(n26) );
  INV2 U68 ( .I(n21), .O(n69) );
  ND3P U69 ( .I1(n43), .I2(n44), .I3(n45), .O(decrypt_shift[4]) );
  INV3 U70 ( .I(n10), .O(n6) );
  INV3 U71 ( .I(n10), .O(n7) );
  BUF2 U72 ( .I(n84), .O(n61) );
  BUF2 U73 ( .I(n10), .O(n83) );
  BUF2 U74 ( .I(n86), .O(n9) );
  BUF2 U75 ( .I(n83), .O(n81) );
  BUF2 U76 ( .I(n86), .O(n10) );
  BUF1 U77 ( .I(n10), .O(n85) );
  BUF2 U78 ( .I(n9), .O(n84) );
  OA12 U79 ( .B1(n63), .B2(n70), .A1(n77), .O(n75) );
  OAI12S U80 ( .B1(n73), .B2(n72), .A1(n4), .O(n77) );
  BUF2 U81 ( .I(n10), .O(n82) );
  OAI12S U83 ( .B1(n70), .B2(n13), .A1(n71), .O(N66) );
  OR3 U84 ( .I1(n72), .I2(n73), .I3(n63), .O(n71) );
  NR2 U85 ( .I1(n22), .I2(n23), .O(n17) );
  INV2 U86 ( .I(n16), .O(n15) );
  INV2 U87 ( .I(state), .O(n86) );
  NR2 U88 ( .I1(n4), .I2(din_valid), .O(stall) );
  OAI112 U89 ( .C1(n51), .C2(n36), .A1(n52), .B1(n35), .O(decrypt_shift[1]) );
  ND2 U90 ( .I1(n51), .I2(n59), .O(n52) );
  NR2P U91 ( .I1(n60), .I2(edr[0]), .O(n51) );
  BUF2 U92 ( .I(n87), .O(round[0]) );
  INV2 U93 ( .I(round[2]), .O(n18) );
  AO22 U94 ( .A1(dout[47]), .A2(n7), .B1(din[46]), .B2(n84), .O(r_din[58]) );
  AO22 U95 ( .A1(dout[61]), .A2(n7), .B1(din[60]), .B2(n83), .O(r_din[48]) );
  AO22 U96 ( .A1(dout[57]), .A2(n5), .B1(din[56]), .B2(n61), .O(r_din[32]) );
  NR2T U97 ( .I1(round[3]), .I2(round[2]), .O(n66) );
  ND2P U98 ( .I1(round[0]), .I2(round[1]), .O(n29) );
  AO22 U99 ( .A1(dout[25]), .A2(n6), .B1(din[24]), .B2(n81), .O(r_din[36]) );
  AO22 U100 ( .A1(dout[9]), .A2(n6), .B1(din[8]), .B2(n81), .O(r_din[38]) );
  AO22 U101 ( .A1(dout[11]), .A2(n6), .B1(din[10]), .B2(n82), .O(r_din[46]) );
  AO22 U102 ( .A1(dout[3]), .A2(n6), .B1(din[2]), .B2(n82), .O(r_din[47]) );
  AO22 U103 ( .A1(dout[15]), .A2(state), .B1(din[14]), .B2(n85), .O(r_din[62])
         );
  AO22 U104 ( .A1(dout[7]), .A2(state), .B1(din[6]), .B2(n85), .O(r_din[63])
         );
  AO22 U105 ( .A1(dout[53]), .A2(n7), .B1(din[52]), .B2(n83), .O(r_din[49]) );
  AO22 U106 ( .A1(dout[13]), .A2(n7), .B1(din[12]), .B2(n83), .O(r_din[54]) );
  AO22 U107 ( .A1(dout[63]), .A2(n7), .B1(din[62]), .B2(n84), .O(r_din[56]) );
  AO22 U108 ( .A1(dout[41]), .A2(n6), .B1(din[40]), .B2(n81), .O(r_din[34]) );
  AO22 U109 ( .A1(dout[33]), .A2(n6), .B1(din[32]), .B2(n81), .O(r_din[35]) );
  AO22 U110 ( .A1(dout[1]), .A2(n6), .B1(din[0]), .B2(n81), .O(r_din[39]) );
  AO22 U111 ( .A1(dout[59]), .A2(n6), .B1(din[58]), .B2(n82), .O(r_din[40]) );
  AO22 U112 ( .A1(dout[51]), .A2(n6), .B1(din[50]), .B2(n82), .O(r_din[41]) );
  AO22 U113 ( .A1(dout[43]), .A2(n6), .B1(din[42]), .B2(n82), .O(r_din[42]) );
  AO22 U114 ( .A1(dout[35]), .A2(n6), .B1(din[34]), .B2(n82), .O(r_din[43]) );
  AO22 U115 ( .A1(dout[19]), .A2(n6), .B1(din[18]), .B2(n82), .O(r_din[45]) );
  AO22 U116 ( .A1(dout[29]), .A2(n7), .B1(din[28]), .B2(n83), .O(r_din[52]) );
  AO22 U117 ( .A1(dout[21]), .A2(n7), .B1(din[20]), .B2(n83), .O(r_din[53]) );
  AO22 U118 ( .A1(dout[55]), .A2(n7), .B1(din[54]), .B2(n84), .O(r_din[57]) );
  AO22 U119 ( .A1(dout[39]), .A2(n7), .B1(din[38]), .B2(n84), .O(r_din[59]) );
  AO22 U120 ( .A1(dout[31]), .A2(n7), .B1(din[30]), .B2(n84), .O(r_din[60]) );
  AO22 U121 ( .A1(dout[23]), .A2(n7), .B1(din[22]), .B2(n84), .O(r_din[61]) );
  AO22 U122 ( .A1(dout[5]), .A2(n7), .B1(din[4]), .B2(n84), .O(r_din[55]) );
  INV2 U123 ( .I(round[1]), .O(n23) );
  AO22 U124 ( .A1(dout[27]), .A2(n6), .B1(din[26]), .B2(n82), .O(r_din[44]) );
  AO22 U125 ( .A1(dout[17]), .A2(n6), .B1(din[16]), .B2(n81), .O(r_din[37]) );
  AO22 U126 ( .A1(dout[45]), .A2(n7), .B1(din[44]), .B2(n83), .O(r_din[50]) );
  AO22 U127 ( .A1(dout[37]), .A2(n7), .B1(din[36]), .B2(n83), .O(r_din[51]) );
  ND2P U128 ( .I1(edr[1]), .I2(edr[0]), .O(n21) );
  MAOI1P U129 ( .A1(n33), .A2(n21), .B1(edr[1]), .B2(n36), .O(n45) );
  ND2P U130 ( .I1(edr[0]), .I2(n60), .O(n13) );
  INV2 U131 ( .I(edr[1]), .O(n60) );
  AO22 U132 ( .A1(dout[34]), .A2(n4), .B1(din[35]), .B2(n8), .O(r_din[11]) );
  AO22 U133 ( .A1(dout[26]), .A2(n4), .B1(din[27]), .B2(n9), .O(r_din[12]) );
  AO22 U134 ( .A1(dout[18]), .A2(n4), .B1(din[19]), .B2(n9), .O(r_din[13]) );
  AO22 U135 ( .A1(dout[2]), .A2(n4), .B1(din[3]), .B2(n9), .O(r_din[15]) );
  AO22 U136 ( .A1(dout[48]), .A2(n5), .B1(din[49]), .B2(n10), .O(r_din[1]) );
  AO22 U137 ( .A1(dout[32]), .A2(n6), .B1(din[33]), .B2(n81), .O(r_din[3]) );
  AO22 U138 ( .A1(dout[16]), .A2(n7), .B1(din[17]), .B2(n84), .O(r_din[5]) );
  AO22 U139 ( .A1(dout[20]), .A2(n5), .B1(din[21]), .B2(n10), .O(r_din[21]) );
  AO22 U140 ( .A1(dout[12]), .A2(n5), .B1(din[13]), .B2(n81), .O(r_din[22]) );
  AO22 U141 ( .A1(dout[4]), .A2(n6), .B1(din[5]), .B2(n10), .O(r_din[23]) );
  AO22 U142 ( .A1(dout[22]), .A2(n5), .B1(din[23]), .B2(n61), .O(r_din[29]) );
  AO22 U143 ( .A1(dout[14]), .A2(n5), .B1(din[15]), .B2(n61), .O(r_din[30]) );
  AO22 U144 ( .A1(n4), .A2(dout[50]), .B1(din[51]), .B2(n10), .O(r_din[9]) );
  AO22 U145 ( .A1(dout[8]), .A2(n4), .B1(din[9]), .B2(n85), .O(r_din[6]) );
  AO22 U146 ( .A1(dout[42]), .A2(n4), .B1(din[43]), .B2(n8), .O(r_din[10]) );
  AO22 U147 ( .A1(dout[10]), .A2(n4), .B1(din[11]), .B2(n9), .O(r_din[14]) );
  AO22 U148 ( .A1(dout[40]), .A2(n5), .B1(din[41]), .B2(n61), .O(r_din[2]) );
  AO22 U149 ( .A1(dout[54]), .A2(n5), .B1(din[55]), .B2(n10), .O(r_din[25]) );
  AO22 U150 ( .A1(dout[49]), .A2(n5), .B1(din[48]), .B2(n61), .O(r_din[33]) );
  AOI13HS U151 ( .B1(n57), .B2(n20), .B3(n74), .A1(n75), .O(N40) );
  ND2 U152 ( .I1(round[3]), .I2(n29), .O(n74) );
  OA222 U153 ( .A1(n21), .A2(round[1]), .B1(n22), .B2(round[3]), .C1(edr[0]), 
        .C2(round[0]), .O(n16) );
  OR2 U154 ( .I1(edr[0]), .I2(edr[1]), .O(n22) );
  ND2 U155 ( .I1(n16), .I2(n78), .O(n72) );
  AO12 U156 ( .B1(round[1]), .B2(round[2]), .A1(n22), .O(n78) );
  NR2 U157 ( .I1(n75), .I2(n76), .O(N39) );
  XOR2 U158 ( .I1(n29), .I2(round[2]), .O(n76) );
  NR2 U159 ( .I1(n2), .I2(n75), .O(N37) );
  BUF1 U160 ( .I(n87), .O(n2) );
  OA112 U161 ( .C1(n79), .C2(n65), .A1(n38), .B1(n22), .O(n73) );
  OA22 U162 ( .A1(edr[0]), .A2(round[1]), .B1(round[0]), .B2(n21), .O(n79) );
  ND3 U163 ( .I1(n21), .I2(n18), .I3(round[1]), .O(n19) );
  OAI12S U164 ( .B1(n11), .B2(n82), .A1(n12), .O(n80) );
  ND3 U165 ( .I1(n13), .I2(n8), .I3(din_valid), .O(n12) );
  AOI112P U166 ( .C1(round[0]), .C2(edr[0]), .A1(n14), .B1(n15), .O(n11) );
  OAI112S U167 ( .C1(n17), .C2(n18), .A1(n19), .B1(n20), .O(n14) );
  INV2 U168 ( .I(din_valid), .O(n70) );
  QDFZRBS dout_valid_reg ( .D(N66), .TD(test_si), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(dout_valid) );
  QDFZRBS state_reg ( .D(n80), .TD(round[3]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(state) );
  QDFZRBS round_reg_0 ( .D(N37), .TD(dout_valid), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(n87) );
  QDFZRBS round_reg_3 ( .D(N40), .TD(round[2]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(round[3]) );
  QDFZRBS round_reg_1 ( .D(N38), .TD(n87), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(round[1]) );
  QDFZRBS round_reg_2 ( .D(N39), .TD(round[1]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(round[2]) );
endmodule


module SNPS_CLOCK_GATE_OBS_des_dat ( TE, net1811, net1816, hclk, test_se, 
        test_si, test_so );
  input TE, net1811, net1816, hclk, test_se, test_si;
  output test_so;
  wire   net1826, net1828, net1830, net1831;

  AN2 main_gate ( .I1(TE), .I2(hclk), .O(net1826) );
  ND2 nand_0_1 ( .I1(net1816), .I2(TE), .O(net1830) );
  ND2 nand_0_0 ( .I1(net1811), .I2(TE), .O(net1828) );
  XOR2 U3 ( .I1(net1830), .I2(net1828), .O(net1831) );
  QDFZS U1 ( .D(net1831), .TD(test_si), .SEL(test_se), .CK(net1826), .Q(
        test_so) );
endmodule


module POWERMODULE_HIGH_des_dat_0_0 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1802;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1802), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1802) );
endmodule


module POWERMODULE_HIGH_des_dat_0_1 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1802;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1802), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1802) );
endmodule


module SNPS_CLOCK_GATE_OBS_des_iv ( TE, net1850, net1855, hclk, test_se, 
        test_si, test_so );
  input TE, net1850, net1855, hclk, test_se, test_si;
  output test_so;
  wire   net1865, net1867, net1869, net1870;

  AN2 main_gate ( .I1(TE), .I2(hclk), .O(net1865) );
  ND2 nand_0_1 ( .I1(net1855), .I2(TE), .O(net1869) );
  ND2 nand_0_0 ( .I1(net1850), .I2(TE), .O(net1867) );
  XOR2 U3 ( .I1(net1869), .I2(net1867), .O(net1870) );
  QDFZS U1 ( .D(net1870), .TD(test_si), .SEL(test_se), .CK(net1865), .Q(
        test_so) );
endmodule


module POWERMODULE_HIGH_des_iv_0_0 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1841;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1841), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1841) );
endmodule


module POWERMODULE_HIGH_des_iv_0_1 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1841;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1841), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1841) );
endmodule


module SNPS_CLOCK_GATE_OBS_des_key ( TE, net1889, net1894, net1899, net1904, 
        net1909, net1914, hclk, test_se, test_si, test_so );
  input TE, net1889, net1894, net1899, net1904, net1909, net1914, hclk,
         test_se, test_si;
  output test_so;
  wire   net1924, net1926, net1928, net1930, net1932, net1934, net1936,
         net1941, n2, n4;

  AN2 main_gate ( .I1(n4), .I2(hclk), .O(net1924) );
  ND2 nand_0_0 ( .I1(net1889), .I2(n4), .O(net1926) );
  ND2 nand_0_2 ( .I1(net1899), .I2(n4), .O(net1930) );
  ND2 nand_0_1 ( .I1(net1894), .I2(n4), .O(net1928) );
  ND2 nand_0_5 ( .I1(net1914), .I2(n4), .O(net1936) );
  ND2 nand_0_4 ( .I1(net1909), .I2(n4), .O(net1934) );
  ND2 nand_0_3 ( .I1(net1904), .I2(n4), .O(net1932) );
  BUF2 U4 ( .I(TE), .O(n4) );
  XOR3 U5 ( .I1(net1936), .I2(net1934), .I3(net1932), .O(n2) );
  XOR4 U6 ( .I1(net1930), .I2(net1928), .I3(n2), .I4(net1926), .O(net1941) );
  QDFZS U1 ( .D(net1941), .TD(test_si), .SEL(test_se), .CK(net1924), .Q(
        test_so) );
endmodule


module POWERMODULE_HIGH_des_key_0_0 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1880;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1880), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1880) );
endmodule


module POWERMODULE_HIGH_des_key_0_1 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1880;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1880), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1880) );
endmodule


module POWERMODULE_HIGH_des_key_0_2 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1880;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1880), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1880) );
endmodule


module POWERMODULE_HIGH_des_key_0_3 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1880;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1880), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1880) );
endmodule


module POWERMODULE_HIGH_des_key_0_4 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1880;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1880), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1880) );
endmodule


module POWERMODULE_HIGH_des_key_0_5 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1880;

  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
  AN2 main_gate ( .I1(net1880), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1880) );
endmodule


module des_spares_0 ( clk, resetn, test_se, test_si, test_so );
  input clk, resetn, test_se, test_si;
  output test_so;
  wire   spare_tie_low, spare_tie_high, spare_na00, spare_nb00, spare_nc00,
         spare_ne00, spare_na01, spare_nb01, spare_nc01, spare_nd01,
         spare_ne01, spare_ng01, spare_na02, spare_nb02, spare_nc02,
         spare_ne02, spare_na03, spare_nb03, spare_nc03, spare_nd03,
         spare_ne03, spare_nf03, spare_ng03, n3;

  TIE0 SPARE_TIEL ( .O(spare_tie_low) );
  TIE1 SPARE_TIEH ( .O(spare_tie_high) );
  NR2T SPARE_UA00 ( .I1(spare_tie_low), .I2(spare_tie_low), .O(spare_na00) );
  INV4 SPARE_UB00 ( .I(spare_na00), .O(spare_nb00) );
  ND2T SPARE_UC00 ( .I1(spare_tie_high), .I2(spare_tie_high), .O(spare_nc00)
         );
  XNR2P SPARE_UE00 ( .I1(spare_nb00), .I2(spare_nc00), .O(spare_ne00) );
  NR2T SPARE_UA01 ( .I1(spare_tie_low), .I2(spare_tie_low), .O(spare_na01) );
  INV4 SPARE_UB01 ( .I(spare_na01), .O(spare_nb01) );
  ND2T SPARE_UC01 ( .I1(spare_tie_high), .I2(spare_tie_high), .O(spare_nc01)
         );
  INV4 SPARE_UD01 ( .I(spare_nc01), .O(spare_nd01) );
  MUX2P SPARE_UE01 ( .A(spare_nb01), .B(spare_nd01), .S(spare_tie_low), .O(
        spare_ne01) );
  NR3T SPARE_UA02 ( .I1(spare_tie_low), .I2(spare_tie_low), .I3(spare_tie_low), 
        .O(spare_na02) );
  INV4 SPARE_UB02 ( .I(spare_na02), .O(spare_nb02) );
  ND3T SPARE_UC02 ( .I1(spare_tie_high), .I2(spare_tie_high), .I3(
        spare_tie_high), .O(spare_nc02) );
  XNR2P SPARE_UE02 ( .I1(spare_nb02), .I2(spare_nc02), .O(spare_ne02) );
  NR3T SPARE_UA03 ( .I1(spare_tie_low), .I2(spare_tie_low), .I3(spare_tie_low), 
        .O(spare_na03) );
  INV4 SPARE_UB03 ( .I(spare_na03), .O(spare_nb03) );
  ND3T SPARE_UC03 ( .I1(spare_tie_high), .I2(spare_tie_high), .I3(
        spare_tie_high), .O(spare_nc03) );
  INV4 SPARE_UD03 ( .I(spare_nc03), .O(spare_nd03) );
  MUX2P SPARE_UE03 ( .A(spare_nb03), .B(spare_nd03), .S(spare_tie_low), .O(
        spare_ne03) );
  DFZRBS SPARE_UF01 ( .D(spare_ne01), .TD(test_si), .SEL(test_se), .CK(clk), 
        .RB(resetn), .Q(n3), .QB(spare_ng01) );
  DFZRBS SPARE_UF03 ( .D(spare_ne03), .TD(n3), .SEL(test_se), .CK(clk), .RB(
        resetn), .Q(spare_nf03), .QB(spare_ng03) );
  QDBHN LOCKUP ( .CKB(clk), .D(spare_nf03), .Q(test_so) );
endmodule


module SNPS_CLOCK_GATE_OBS_des ( TE, net1749, hclk, test_se, test_si, test_so
 );
  input TE, net1749, hclk, test_se, test_si;
  output test_so;
  wire   net1759, net1761;

  AN2 main_gate ( .I1(TE), .I2(hclk), .O(net1759) );
  ND2 nand_0_0 ( .I1(net1749), .I2(TE), .O(net1761) );
  QDFZS U1 ( .D(net1761), .TD(test_si), .SEL(test_se), .CK(net1759), .Q(
        test_so) );
endmodule


module POWERMODULE_HIGH_des_0 ( CLK, EN, ENCLK, TE, ENOBS );
  input CLK, EN, TE;
  output ENCLK, ENOBS;
  wire   net1740;

  AN2 main_gate ( .I1(net1740), .I2(CLK), .O(ENCLK) );
  OR2 U2 ( .I1(TE), .I2(ENOBS), .O(net1740) );
  QDBHN latch ( .CKB(CLK), .D(EN), .Q(ENOBS) );
endmodule


module des_cop ( hclk, POR, hresetn, encrypt_whole, dt_sel, key23_sel, edr, 
        mode_sel, iv_sel, iv, key1, key2, key3, din, din_valid_whole, dout, 
        dout_valid, test_mode, test_se, test_si, test_so );
  input [1:0] edr;
  input [63:0] iv;
  input [63:0] key1;
  input [63:0] key2;
  input [63:0] key3;
  input [63:0] din;
  output [63:0] dout;
  input hclk, POR, hresetn, encrypt_whole, dt_sel, key23_sel, mode_sel, iv_sel,
         din_valid_whole, test_mode, test_se, test_si;
  output dout_valid, test_so;
  wire   encrypt_eins, din_valid_eins, dout_valid_eins, N31, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n27,
         n28, n29, n30, n31, n32, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n26, n33, n34, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, flag_0_;
  wire   [63:0] key_eins;
  wire   [63:0] din_eins;
  wire   [3:0] round;
  wire   [63:0] dout_eins;

  tiny_des des_unit ( .hclk(hclk), .POR(POR), .hresetn(hresetn), .encrypt(
        encrypt_eins), .edr(edr), .key_in(key_eins), .din(din_eins), 
        .din_valid(din_valid_eins), .round(round), .dout(dout_eins), 
        .dout_valid(dout_valid_eins), .test_mode(test_mode), .test_se(test_se), 
        .test_si(test_si) );
  OR2P U3 ( .I1(n295), .I2(flag_0_), .O(n1) );
  ND2 U4 ( .I1(flag_0_), .I2(n295), .O(n29) );
  ND2P U5 ( .I1(n297), .I2(n31), .O(n168) );
  BUF1 U6 ( .I(n10), .O(n343) );
  BUF2 U7 ( .I(n10), .O(n335) );
  BUF2 U8 ( .I(n10), .O(n341) );
  BUF2 U9 ( .I(n10), .O(n336) );
  BUF2 U10 ( .I(n10), .O(n334) );
  BUF2 U11 ( .I(n10), .O(n342) );
  BUF2 U12 ( .I(n10), .O(n340) );
  BUF2 U13 ( .I(n10), .O(n339) );
  BUF2 U14 ( .I(n10), .O(n338) );
  BUF2 U15 ( .I(n10), .O(n337) );
  AO222 U16 ( .A1(key3[0]), .A2(n333), .B1(key1[0]), .B2(n329), .C1(key2[0]), 
        .C2(n325), .O(key_eins[0]) );
  AO222 U17 ( .A1(key3[16]), .A2(n333), .B1(key1[16]), .B2(n329), .C1(key2[16]), .C2(n325), .O(key_eins[16]) );
  AO222 U18 ( .A1(key3[24]), .A2(n332), .B1(key1[24]), .B2(n328), .C1(key2[24]), .C2(n324), .O(key_eins[24]) );
  AO222 U19 ( .A1(key3[32]), .A2(n332), .B1(key1[32]), .B2(n328), .C1(key2[32]), .C2(n324), .O(key_eins[32]) );
  AO222 U20 ( .A1(key3[40]), .A2(n331), .B1(key1[40]), .B2(n327), .C1(key2[40]), .C2(n323), .O(key_eins[40]) );
  AO222 U21 ( .A1(key3[48]), .A2(n331), .B1(key1[48]), .B2(n327), .C1(key2[48]), .C2(n323), .O(key_eins[48]) );
  AO222 U22 ( .A1(key3[56]), .A2(n330), .B1(key1[56]), .B2(n326), .C1(key2[56]), .C2(n322), .O(key_eins[56]) );
  AO222 U23 ( .A1(key3[8]), .A2(n330), .B1(key1[8]), .B2(n326), .C1(key2[8]), 
        .C2(n322), .O(key_eins[8]) );
  INV3 U24 ( .I(n31), .O(n10) );
  BUF2 U25 ( .I(n25), .O(n329) );
  BUF2 U26 ( .I(n25), .O(n328) );
  BUF2 U27 ( .I(n25), .O(n327) );
  BUF2 U28 ( .I(n25), .O(n326) );
  INV3 U29 ( .I(n1), .O(n325) );
  INV3 U30 ( .I(n1), .O(n323) );
  INV3 U31 ( .I(n1), .O(n322) );
  INV3 U32 ( .I(n1), .O(n324) );
  BUF2 U33 ( .I(n24), .O(n333) );
  BUF2 U34 ( .I(n24), .O(n332) );
  BUF2 U35 ( .I(n24), .O(n331) );
  BUF2 U36 ( .I(n24), .O(n330) );
  BUF2 U37 ( .I(n167), .O(n306) );
  BUF2 U38 ( .I(n167), .O(n308) );
  BUF2 U39 ( .I(n167), .O(n307) );
  BUF2 U40 ( .I(n167), .O(n309) );
  ND2P U41 ( .I1(n16), .I2(n295), .O(n22) );
  OAI112 U42 ( .C1(n343), .C2(n27), .A1(n28), .B1(n22), .O(n25) );
  OR2B1 U43 ( .I1(n29), .B1(n30), .O(n28) );
  NR2P U44 ( .I1(n295), .I2(n16), .O(n31) );
  MOAI1P U45 ( .A1(n30), .A2(n29), .B1(n31), .B2(n27), .O(n24) );
  BUF2 U46 ( .I(n166), .O(n310) );
  BUF1 U47 ( .I(n168), .O(n9) );
  BUF1 U48 ( .I(n168), .O(n3) );
  BUF1 U49 ( .I(n168), .O(n26) );
  BUF1 U50 ( .I(n168), .O(n33) );
  BUF1 U51 ( .I(n168), .O(n2) );
  ND3P U52 ( .I1(n29), .I2(n22), .I3(n1), .O(n167) );
  BUF2 U53 ( .I(n166), .O(n311) );
  BUF2 U54 ( .I(n166), .O(n312) );
  BUF2 U55 ( .I(n166), .O(n313) );
  BUF1 U56 ( .I(n168), .O(n6) );
  BUF1 U57 ( .I(n168), .O(n4) );
  BUF1 U58 ( .I(n168), .O(n5) );
  BUF1 U59 ( .I(n168), .O(n7) );
  BUF1 U60 ( .I(n168), .O(n8) );
  BUF1 U61 ( .I(n168), .O(n34) );
  ND3 U62 ( .I1(n18), .I2(n19), .I3(n20), .O(n14) );
  AN3 U63 ( .I1(n21), .I2(n22), .I3(n23), .O(n20) );
  ND2 U64 ( .I1(n303), .I2(n302), .O(n300) );
  BUF2 U65 ( .I(n36), .O(n317) );
  BUF2 U66 ( .I(n36), .O(n316) );
  BUF2 U67 ( .I(n36), .O(n315) );
  BUF2 U68 ( .I(n36), .O(n314) );
  BUF2 U69 ( .I(n36), .O(n321) );
  BUF2 U70 ( .I(n36), .O(n320) );
  BUF2 U71 ( .I(n36), .O(n319) );
  BUF2 U72 ( .I(n36), .O(n318) );
  INV2 U73 ( .I(test_so), .O(n295) );
  AN2B1 U74 ( .I1(dout_valid_eins), .B1(n22), .O(dout_valid) );
  INV2 U75 ( .I(flag_0_), .O(n16) );
  AO222 U76 ( .A1(key3[37]), .A2(n332), .B1(key1[37]), .B2(n328), .C1(key2[37]), .C2(n324), .O(key_eins[37]) );
  AO222 U77 ( .A1(key3[4]), .A2(n331), .B1(key1[4]), .B2(n327), .C1(key2[4]), 
        .C2(n323), .O(key_eins[4]) );
  AO222 U78 ( .A1(key3[7]), .A2(n330), .B1(key1[7]), .B2(n326), .C1(key2[7]), 
        .C2(n322), .O(key_eins[7]) );
  AO222 U79 ( .A1(key3[6]), .A2(n330), .B1(key1[6]), .B2(n326), .C1(key2[6]), 
        .C2(n322), .O(key_eins[6]) );
  AO222 U80 ( .A1(key3[38]), .A2(n332), .B1(key1[38]), .B2(n328), .C1(key2[38]), .C2(n324), .O(key_eins[38]) );
  AO222 U81 ( .A1(key3[29]), .A2(n332), .B1(key1[29]), .B2(n328), .C1(key2[29]), .C2(n324), .O(key_eins[29]) );
  AO222 U82 ( .A1(key3[61]), .A2(n330), .B1(key1[61]), .B2(n326), .C1(key2[61]), .C2(n322), .O(key_eins[61]) );
  AO222 U83 ( .A1(key3[31]), .A2(n332), .B1(key1[31]), .B2(n328), .C1(key2[31]), .C2(n324), .O(key_eins[31]) );
  AO222 U84 ( .A1(key3[30]), .A2(n332), .B1(key1[30]), .B2(n328), .C1(key2[30]), .C2(n324), .O(key_eins[30]) );
  AO222 U85 ( .A1(key3[45]), .A2(n331), .B1(key1[45]), .B2(n327), .C1(key2[45]), .C2(n323), .O(key_eins[45]) );
  AO222 U86 ( .A1(key3[47]), .A2(n331), .B1(key1[47]), .B2(n327), .C1(key2[47]), .C2(n323), .O(key_eins[47]) );
  AO222 U87 ( .A1(key3[15]), .A2(n333), .B1(key1[15]), .B2(n329), .C1(key2[15]), .C2(n325), .O(key_eins[15]) );
  AO222 U88 ( .A1(key3[12]), .A2(n333), .B1(key1[12]), .B2(n329), .C1(key2[12]), .C2(n325), .O(key_eins[12]) );
  AO222 U89 ( .A1(key3[46]), .A2(n331), .B1(key1[46]), .B2(n327), .C1(key2[46]), .C2(n323), .O(key_eins[46]) );
  AO222 U90 ( .A1(key3[5]), .A2(n330), .B1(key1[5]), .B2(n326), .C1(key2[5]), 
        .C2(n322), .O(key_eins[5]) );
  AO222 U91 ( .A1(key3[62]), .A2(n330), .B1(key1[62]), .B2(n326), .C1(key2[62]), .C2(n322), .O(key_eins[62]) );
  AO222 U92 ( .A1(key3[21]), .A2(n333), .B1(key1[21]), .B2(n329), .C1(key2[21]), .C2(n325), .O(key_eins[21]) );
  AO222 U93 ( .A1(key3[20]), .A2(n333), .B1(key1[20]), .B2(n329), .C1(key2[20]), .C2(n325), .O(key_eins[20]) );
  AO222 U94 ( .A1(key3[54]), .A2(n330), .B1(key1[54]), .B2(n326), .C1(key2[54]), .C2(n322), .O(key_eins[54]) );
  AO222 U95 ( .A1(key3[13]), .A2(n333), .B1(key1[13]), .B2(n329), .C1(key2[13]), .C2(n325), .O(key_eins[13]) );
  AO222 U96 ( .A1(key3[53]), .A2(n330), .B1(key1[53]), .B2(n326), .C1(key2[53]), .C2(n322), .O(key_eins[53]) );
  AO222 U97 ( .A1(key3[55]), .A2(n330), .B1(key1[55]), .B2(n326), .C1(key2[55]), .C2(n322), .O(key_eins[55]) );
  AO222 U98 ( .A1(key3[63]), .A2(n330), .B1(key1[63]), .B2(n326), .C1(key2[63]), .C2(n322), .O(key_eins[63]) );
  AO222 U99 ( .A1(key3[28]), .A2(n332), .B1(key1[28]), .B2(n328), .C1(key2[28]), .C2(n324), .O(key_eins[28]) );
  AO222 U100 ( .A1(key3[22]), .A2(n333), .B1(key1[22]), .B2(n329), .C1(
        key2[22]), .C2(n325), .O(key_eins[22]) );
  AN3 U101 ( .I1(mode_sel), .I2(iv_sel), .I3(n296), .O(n166) );
  NR2 U102 ( .I1(encrypt_whole), .I2(n343), .O(n296) );
  AO222 U103 ( .A1(key3[44]), .A2(n331), .B1(key1[44]), .B2(n327), .C1(
        key2[44]), .C2(n323), .O(key_eins[44]) );
  AO222 U104 ( .A1(key3[42]), .A2(n331), .B1(key1[42]), .B2(n327), .C1(
        key2[42]), .C2(n323), .O(key_eins[42]) );
  AO222 U105 ( .A1(key3[41]), .A2(n331), .B1(key1[41]), .B2(n327), .C1(
        key2[41]), .C2(n323), .O(key_eins[41]) );
  AO222 U106 ( .A1(key3[25]), .A2(n332), .B1(key1[25]), .B2(n328), .C1(
        key2[25]), .C2(n324), .O(key_eins[25]) );
  AO222 U107 ( .A1(key3[59]), .A2(n330), .B1(key1[59]), .B2(n326), .C1(
        key2[59]), .C2(n322), .O(key_eins[59]) );
  AO222 U108 ( .A1(key3[60]), .A2(n330), .B1(key1[60]), .B2(n326), .C1(
        key2[60]), .C2(n322), .O(key_eins[60]) );
  AO222 U109 ( .A1(key3[57]), .A2(n330), .B1(key1[57]), .B2(n326), .C1(
        key2[57]), .C2(n322), .O(key_eins[57]) );
  AO222 U110 ( .A1(key3[58]), .A2(n330), .B1(key1[58]), .B2(n326), .C1(
        key2[58]), .C2(n322), .O(key_eins[58]) );
  AO222 U111 ( .A1(key3[26]), .A2(n332), .B1(key1[26]), .B2(n328), .C1(
        key2[26]), .C2(n324), .O(key_eins[26]) );
  AO222 U112 ( .A1(key3[27]), .A2(n332), .B1(key1[27]), .B2(n328), .C1(
        key2[27]), .C2(n324), .O(key_eins[27]) );
  AO222 U113 ( .A1(key3[17]), .A2(n333), .B1(key1[17]), .B2(n329), .C1(
        key2[17]), .C2(n325), .O(key_eins[17]) );
  AO222 U114 ( .A1(key3[50]), .A2(n331), .B1(key1[50]), .B2(n327), .C1(
        key2[50]), .C2(n323), .O(key_eins[50]) );
  AO222 U115 ( .A1(key3[18]), .A2(n333), .B1(key1[18]), .B2(n329), .C1(
        key2[18]), .C2(n325), .O(key_eins[18]) );
  AO222 U116 ( .A1(key3[36]), .A2(n332), .B1(key1[36]), .B2(n328), .C1(
        key2[36]), .C2(n324), .O(key_eins[36]) );
  AO222 U117 ( .A1(key3[1]), .A2(n333), .B1(key1[1]), .B2(n329), .C1(key2[1]), 
        .C2(n325), .O(key_eins[1]) );
  AO222 U118 ( .A1(key3[2]), .A2(n332), .B1(key1[2]), .B2(n328), .C1(key2[2]), 
        .C2(n324), .O(key_eins[2]) );
  AO222 U119 ( .A1(key3[39]), .A2(n331), .B1(key1[39]), .B2(n327), .C1(
        key2[39]), .C2(n323), .O(key_eins[39]) );
  AO222 U120 ( .A1(key3[14]), .A2(n333), .B1(key1[14]), .B2(n329), .C1(
        key2[14]), .C2(n325), .O(key_eins[14]) );
  AO222 U121 ( .A1(key3[23]), .A2(n333), .B1(key1[23]), .B2(n329), .C1(
        key2[23]), .C2(n325), .O(key_eins[23]) );
  AO222 U122 ( .A1(key3[33]), .A2(n332), .B1(key1[33]), .B2(n328), .C1(
        key2[33]), .C2(n324), .O(key_eins[33]) );
  AO222 U123 ( .A1(key3[51]), .A2(n331), .B1(key1[51]), .B2(n327), .C1(
        key2[51]), .C2(n323), .O(key_eins[51]) );
  AO222 U124 ( .A1(key3[52]), .A2(n331), .B1(key1[52]), .B2(n327), .C1(
        key2[52]), .C2(n323), .O(key_eins[52]) );
  AO222 U125 ( .A1(key3[9]), .A2(n330), .B1(key1[9]), .B2(n326), .C1(key2[9]), 
        .C2(n322), .O(key_eins[9]) );
  AO222 U126 ( .A1(key3[43]), .A2(n331), .B1(key1[43]), .B2(n327), .C1(
        key2[43]), .C2(n323), .O(key_eins[43]) );
  AO222 U127 ( .A1(key3[49]), .A2(n331), .B1(key1[49]), .B2(n327), .C1(
        key2[49]), .C2(n323), .O(key_eins[49]) );
  AO222 U128 ( .A1(key3[3]), .A2(n331), .B1(key1[3]), .B2(n327), .C1(key2[3]), 
        .C2(n323), .O(key_eins[3]) );
  AO222 U129 ( .A1(key3[34]), .A2(n332), .B1(key1[34]), .B2(n328), .C1(
        key2[34]), .C2(n324), .O(key_eins[34]) );
  AO222 U130 ( .A1(key3[10]), .A2(n333), .B1(key1[10]), .B2(n329), .C1(
        key2[10]), .C2(n325), .O(key_eins[10]) );
  AO222 U131 ( .A1(key3[35]), .A2(n332), .B1(key1[35]), .B2(n328), .C1(
        key2[35]), .C2(n324), .O(key_eins[35]) );
  AO222 U132 ( .A1(key3[19]), .A2(n333), .B1(key1[19]), .B2(n329), .C1(
        key2[19]), .C2(n325), .O(key_eins[19]) );
  AO222 U133 ( .A1(key3[11]), .A2(n333), .B1(key1[11]), .B2(n329), .C1(
        key2[11]), .C2(n325), .O(key_eins[11]) );
  AN3 U134 ( .I1(key23_sel), .I2(dt_sel), .I3(encrypt_whole), .O(n27) );
  INV2 U135 ( .I(encrypt_whole), .O(n32) );
  ND2 U136 ( .I1(key23_sel), .I2(n32), .O(n30) );
  AO222 U137 ( .A1(din[63]), .A2(n175), .B1(n176), .B2(n310), .C1(
        dout_eins[63]), .C2(n306), .O(din_eins[63]) );
  NR2 U138 ( .I1(din[63]), .I2(n45), .O(n176) );
  OAI12S U139 ( .B1(iv[63]), .B2(n342), .A1(n2), .O(n175) );
  AO222 U140 ( .A1(din[25]), .A2(n259), .B1(n260), .B2(n312), .C1(
        dout_eins[25]), .C2(n308), .O(din_eins[25]) );
  NR2 U141 ( .I1(din[25]), .I2(n129), .O(n260) );
  OAI12S U142 ( .B1(iv[25]), .B2(n336), .A1(n9), .O(n259) );
  AO222 U143 ( .A1(din[37]), .A2(n233), .B1(n234), .B2(n312), .C1(
        dout_eins[37]), .C2(n308), .O(din_eins[37]) );
  NR2 U144 ( .I1(din[37]), .I2(n103), .O(n234) );
  OAI12S U145 ( .B1(iv[37]), .B2(n338), .A1(n7), .O(n233) );
  AO222 U146 ( .A1(din[29]), .A2(n251), .B1(n252), .B2(n312), .C1(
        dout_eins[29]), .C2(n308), .O(din_eins[29]) );
  NR2 U147 ( .I1(din[29]), .I2(n121), .O(n252) );
  OAI12S U148 ( .B1(iv[29]), .B2(n336), .A1(n9), .O(n251) );
  AO222 U149 ( .A1(din[39]), .A2(n229), .B1(n230), .B2(n311), .C1(
        dout_eins[39]), .C2(n307), .O(din_eins[39]) );
  NR2 U150 ( .I1(din[39]), .I2(n99), .O(n230) );
  OAI12S U151 ( .B1(iv[39]), .B2(n338), .A1(n7), .O(n229) );
  ND3 U152 ( .I1(iv_sel), .I2(n32), .I3(mode_sel), .O(n297) );
  AO222 U153 ( .A1(din[57]), .A2(n189), .B1(n190), .B2(n310), .C1(
        dout_eins[57]), .C2(n306), .O(din_eins[57]) );
  NR2 U154 ( .I1(din[57]), .I2(n59), .O(n190) );
  OAI12S U155 ( .B1(iv[57]), .B2(n341), .A1(n3), .O(n189) );
  AO222 U156 ( .A1(din[31]), .A2(n245), .B1(n246), .B2(n312), .C1(
        dout_eins[31]), .C2(n308), .O(din_eins[31]) );
  NR2 U157 ( .I1(din[31]), .I2(n115), .O(n246) );
  OAI12S U158 ( .B1(iv[31]), .B2(n337), .A1(n8), .O(n245) );
  AO222 U159 ( .A1(din[7]), .A2(n171), .B1(n172), .B2(n310), .C1(dout_eins[7]), 
        .C2(n306), .O(din_eins[7]) );
  NR2 U160 ( .I1(din[7]), .I2(n41), .O(n172) );
  OAI12S U161 ( .B1(iv[7]), .B2(n342), .A1(n2), .O(n171) );
  AO222 U162 ( .A1(din[1]), .A2(n271), .B1(n272), .B2(n313), .C1(dout_eins[1]), 
        .C2(n309), .O(din_eins[1]) );
  NR2 U163 ( .I1(din[1]), .I2(n141), .O(n272) );
  OAI12S U164 ( .B1(iv[1]), .B2(n335), .A1(n26), .O(n271) );
  AO222 U165 ( .A1(din[59]), .A2(n185), .B1(n186), .B2(n310), .C1(
        dout_eins[59]), .C2(n306), .O(din_eins[59]) );
  NR2 U166 ( .I1(din[59]), .I2(n55), .O(n186) );
  OAI12S U167 ( .B1(iv[59]), .B2(n341), .A1(n3), .O(n185) );
  AO222 U168 ( .A1(din[53]), .A2(n197), .B1(n198), .B2(n310), .C1(
        dout_eins[53]), .C2(n306), .O(din_eins[53]) );
  NR2 U169 ( .I1(din[53]), .I2(n67), .O(n198) );
  OAI12S U170 ( .B1(iv[53]), .B2(n340), .A1(n4), .O(n197) );
  AO222 U171 ( .A1(din[61]), .A2(n179), .B1(n180), .B2(n310), .C1(
        dout_eins[61]), .C2(n306), .O(din_eins[61]) );
  NR2 U172 ( .I1(din[61]), .I2(n49), .O(n180) );
  OAI12S U173 ( .B1(iv[61]), .B2(n342), .A1(n3), .O(n179) );
  AO222 U174 ( .A1(din[47]), .A2(n211), .B1(n212), .B2(n311), .C1(
        dout_eins[47]), .C2(n307), .O(din_eins[47]) );
  NR2 U175 ( .I1(din[47]), .I2(n81), .O(n212) );
  OAI12S U176 ( .B1(iv[47]), .B2(n339), .A1(n5), .O(n211) );
  AO222 U177 ( .A1(din[35]), .A2(n237), .B1(n238), .B2(n312), .C1(
        dout_eins[35]), .C2(n308), .O(din_eins[35]) );
  NR2 U178 ( .I1(din[35]), .I2(n107), .O(n238) );
  OAI12S U179 ( .B1(iv[35]), .B2(n337), .A1(n7), .O(n237) );
  AO222 U180 ( .A1(din[27]), .A2(n255), .B1(n256), .B2(n312), .C1(
        dout_eins[27]), .C2(n308), .O(din_eins[27]) );
  NR2 U181 ( .I1(din[27]), .I2(n125), .O(n256) );
  OAI12S U182 ( .B1(iv[27]), .B2(n336), .A1(n9), .O(n255) );
  AO222 U183 ( .A1(din[19]), .A2(n273), .B1(n274), .B2(n313), .C1(
        dout_eins[19]), .C2(n309), .O(din_eins[19]) );
  NR2 U184 ( .I1(din[19]), .I2(n143), .O(n274) );
  OAI12S U185 ( .B1(iv[19]), .B2(n335), .A1(n26), .O(n273) );
  AO222 U186 ( .A1(din[3]), .A2(n227), .B1(n228), .B2(n311), .C1(dout_eins[3]), 
        .C2(n307), .O(din_eins[3]) );
  NR2 U187 ( .I1(din[3]), .I2(n97), .O(n228) );
  OAI12S U188 ( .B1(iv[3]), .B2(n338), .A1(n7), .O(n227) );
  AO222 U189 ( .A1(din[49]), .A2(n207), .B1(n208), .B2(n311), .C1(
        dout_eins[49]), .C2(n307), .O(din_eins[49]) );
  NR2 U190 ( .I1(din[49]), .I2(n77), .O(n208) );
  OAI12S U191 ( .B1(iv[49]), .B2(n340), .A1(n5), .O(n207) );
  AO222 U192 ( .A1(din[33]), .A2(n241), .B1(n242), .B2(n312), .C1(
        dout_eins[33]), .C2(n308), .O(din_eins[33]) );
  NR2 U193 ( .I1(din[33]), .I2(n111), .O(n242) );
  OAI12S U194 ( .B1(iv[33]), .B2(n337), .A1(n8), .O(n241) );
  AO222 U195 ( .A1(din[17]), .A2(n277), .B1(n278), .B2(n313), .C1(
        dout_eins[17]), .C2(n309), .O(din_eins[17]) );
  NR2 U196 ( .I1(din[17]), .I2(n147), .O(n278) );
  OAI12S U197 ( .B1(iv[17]), .B2(n335), .A1(n33), .O(n277) );
  AO222 U198 ( .A1(din[21]), .A2(n267), .B1(n268), .B2(n313), .C1(
        dout_eins[21]), .C2(n309), .O(din_eins[21]) );
  NR2 U199 ( .I1(din[21]), .I2(n137), .O(n268) );
  OAI12S U200 ( .B1(iv[21]), .B2(n335), .A1(n26), .O(n267) );
  AO222 U201 ( .A1(din[13]), .A2(n285), .B1(n286), .B2(n313), .C1(
        dout_eins[13]), .C2(n309), .O(din_eins[13]) );
  NR2 U202 ( .I1(din[13]), .I2(n155), .O(n286) );
  OAI12S U203 ( .B1(iv[13]), .B2(n334), .A1(n33), .O(n285) );
  AO222 U204 ( .A1(din[5]), .A2(n183), .B1(n184), .B2(n310), .C1(dout_eins[5]), 
        .C2(n306), .O(din_eins[5]) );
  NR2 U205 ( .I1(din[5]), .I2(n53), .O(n184) );
  OAI12S U206 ( .B1(iv[5]), .B2(n341), .A1(n3), .O(n183) );
  AO222 U207 ( .A1(din[23]), .A2(n263), .B1(n264), .B2(n313), .C1(
        dout_eins[23]), .C2(n309), .O(din_eins[23]) );
  NR2 U208 ( .I1(din[23]), .I2(n133), .O(n264) );
  OAI12S U209 ( .B1(iv[23]), .B2(n336), .A1(n26), .O(n263) );
  AO222 U210 ( .A1(din[15]), .A2(n281), .B1(n282), .B2(n313), .C1(
        dout_eins[15]), .C2(n309), .O(din_eins[15]) );
  NR2 U211 ( .I1(din[15]), .I2(n151), .O(n282) );
  OAI12S U212 ( .B1(iv[15]), .B2(n334), .A1(n33), .O(n281) );
  AO222 U213 ( .A1(din[51]), .A2(n201), .B1(n202), .B2(n311), .C1(
        dout_eins[51]), .C2(n307), .O(din_eins[51]) );
  NR2 U214 ( .I1(din[51]), .I2(n71), .O(n202) );
  OAI12S U215 ( .B1(iv[51]), .B2(n340), .A1(n4), .O(n201) );
  AO222 U216 ( .A1(din[9]), .A2(n164), .B1(n165), .B2(n310), .C1(dout_eins[9]), 
        .C2(n306), .O(din_eins[9]) );
  NR2 U217 ( .I1(din[9]), .I2(n37), .O(n165) );
  OAI12S U218 ( .B1(iv[9]), .B2(n343), .A1(n2), .O(n164) );
  AO222 U219 ( .A1(din[43]), .A2(n219), .B1(n220), .B2(n311), .C1(
        dout_eins[43]), .C2(n307), .O(din_eins[43]) );
  NR2 U220 ( .I1(din[43]), .I2(n89), .O(n220) );
  OAI12S U221 ( .B1(iv[43]), .B2(n339), .A1(n6), .O(n219) );
  AO222 U222 ( .A1(din[11]), .A2(n289), .B1(n290), .B2(n313), .C1(
        dout_eins[11]), .C2(n309), .O(din_eins[11]) );
  NR2 U223 ( .I1(din[11]), .I2(n159), .O(n290) );
  OAI12S U224 ( .B1(iv[11]), .B2(n334), .A1(n34), .O(n289) );
  AO222 U225 ( .A1(din[41]), .A2(n223), .B1(n224), .B2(n311), .C1(
        dout_eins[41]), .C2(n307), .O(din_eins[41]) );
  NR2 U226 ( .I1(din[41]), .I2(n93), .O(n224) );
  OAI12S U227 ( .B1(iv[41]), .B2(n339), .A1(n6), .O(n223) );
  AO222 U228 ( .A1(din[45]), .A2(n215), .B1(n216), .B2(n311), .C1(
        dout_eins[45]), .C2(n307), .O(din_eins[45]) );
  NR2 U229 ( .I1(din[45]), .I2(n85), .O(n216) );
  OAI12S U230 ( .B1(iv[45]), .B2(n339), .A1(n6), .O(n215) );
  AO222 U231 ( .A1(din[55]), .A2(n193), .B1(n194), .B2(n310), .C1(
        dout_eins[55]), .C2(n306), .O(din_eins[55]) );
  NR2 U232 ( .I1(din[55]), .I2(n63), .O(n194) );
  OAI12S U233 ( .B1(iv[55]), .B2(n341), .A1(n4), .O(n193) );
  INV2 U234 ( .I(iv[63]), .O(n45) );
  INV2 U235 ( .I(iv[33]), .O(n111) );
  INV2 U236 ( .I(iv[35]), .O(n107) );
  INV2 U237 ( .I(iv[37]), .O(n103) );
  INV2 U238 ( .I(iv[39]), .O(n99) );
  INV2 U239 ( .I(iv[47]), .O(n81) );
  INV2 U240 ( .I(iv[49]), .O(n77) );
  INV2 U241 ( .I(iv[51]), .O(n71) );
  INV2 U242 ( .I(iv[53]), .O(n67) );
  INV2 U243 ( .I(iv[57]), .O(n59) );
  INV2 U244 ( .I(iv[59]), .O(n55) );
  INV2 U245 ( .I(iv[61]), .O(n49) );
  INV2 U246 ( .I(iv[1]), .O(n141) );
  INV2 U247 ( .I(iv[3]), .O(n97) );
  INV2 U248 ( .I(iv[5]), .O(n53) );
  INV2 U249 ( .I(iv[7]), .O(n41) );
  INV2 U250 ( .I(iv[9]), .O(n37) );
  INV2 U251 ( .I(iv[11]), .O(n159) );
  INV2 U252 ( .I(iv[13]), .O(n155) );
  INV2 U253 ( .I(iv[17]), .O(n147) );
  INV2 U254 ( .I(iv[19]), .O(n143) );
  INV2 U255 ( .I(iv[21]), .O(n137) );
  INV2 U256 ( .I(iv[23]), .O(n133) );
  INV2 U257 ( .I(iv[25]), .O(n129) );
  INV2 U258 ( .I(iv[27]), .O(n125) );
  INV2 U259 ( .I(iv[29]), .O(n121) );
  INV2 U260 ( .I(iv[31]), .O(n115) );
  INV2 U261 ( .I(iv[41]), .O(n93) );
  INV2 U262 ( .I(iv[43]), .O(n89) );
  INV2 U263 ( .I(iv[45]), .O(n85) );
  INV2 U264 ( .I(iv[55]), .O(n63) );
  INV2 U265 ( .I(iv[15]), .O(n151) );
  AO222 U266 ( .A1(din[48]), .A2(n209), .B1(n210), .B2(n311), .C1(
        dout_eins[48]), .C2(n307), .O(din_eins[48]) );
  NR2 U267 ( .I1(din[48]), .I2(n79), .O(n210) );
  OAI12S U268 ( .B1(iv[48]), .B2(n340), .A1(n5), .O(n209) );
  AO222 U269 ( .A1(din[56]), .A2(n191), .B1(n192), .B2(n310), .C1(
        dout_eins[56]), .C2(n306), .O(din_eins[56]) );
  NR2 U270 ( .I1(din[56]), .I2(n61), .O(n192) );
  OAI12S U271 ( .B1(iv[56]), .B2(n341), .A1(n4), .O(n191) );
  AO222 U272 ( .A1(din[40]), .A2(n225), .B1(n226), .B2(n311), .C1(
        dout_eins[40]), .C2(n307), .O(din_eins[40]) );
  NR2 U273 ( .I1(din[40]), .I2(n95), .O(n226) );
  OAI12S U274 ( .B1(iv[40]), .B2(n338), .A1(n6), .O(n225) );
  AO222 U275 ( .A1(din[32]), .A2(n243), .B1(n244), .B2(n312), .C1(
        dout_eins[32]), .C2(n308), .O(din_eins[32]) );
  NR2 U276 ( .I1(din[32]), .I2(n113), .O(n244) );
  OAI12S U277 ( .B1(iv[32]), .B2(n337), .A1(n8), .O(n243) );
  AO222 U278 ( .A1(din[24]), .A2(n261), .B1(n262), .B2(n312), .C1(
        dout_eins[24]), .C2(n308), .O(din_eins[24]) );
  NR2 U279 ( .I1(din[24]), .I2(n131), .O(n262) );
  OAI12S U280 ( .B1(iv[24]), .B2(n336), .A1(n9), .O(n261) );
  AO222 U281 ( .A1(din[16]), .A2(n279), .B1(n280), .B2(n313), .C1(
        dout_eins[16]), .C2(n309), .O(din_eins[16]) );
  NR2 U282 ( .I1(din[16]), .I2(n149), .O(n280) );
  OAI12S U283 ( .B1(iv[16]), .B2(n334), .A1(n33), .O(n279) );
  AO222 U284 ( .A1(din[8]), .A2(n169), .B1(n170), .B2(n310), .C1(dout_eins[8]), 
        .C2(n306), .O(din_eins[8]) );
  NR2 U285 ( .I1(din[8]), .I2(n39), .O(n170) );
  OAI12S U286 ( .B1(iv[8]), .B2(n342), .A1(n2), .O(n169) );
  AO222 U287 ( .A1(din[0]), .A2(n293), .B1(n294), .B2(n313), .C1(dout_eins[0]), 
        .C2(n309), .O(din_eins[0]) );
  NR2 U288 ( .I1(din[0]), .I2(n163), .O(n294) );
  OAI12S U289 ( .B1(iv[0]), .B2(n338), .A1(n34), .O(n293) );
  AO222 U290 ( .A1(din[58]), .A2(n187), .B1(n188), .B2(n310), .C1(
        dout_eins[58]), .C2(n306), .O(din_eins[58]) );
  NR2 U291 ( .I1(din[58]), .I2(n57), .O(n188) );
  OAI12S U292 ( .B1(iv[58]), .B2(n341), .A1(n3), .O(n187) );
  AO222 U293 ( .A1(din[50]), .A2(n203), .B1(n204), .B2(n311), .C1(
        dout_eins[50]), .C2(n307), .O(din_eins[50]) );
  NR2 U294 ( .I1(din[50]), .I2(n73), .O(n204) );
  OAI12S U295 ( .B1(iv[50]), .B2(n340), .A1(n5), .O(n203) );
  AO222 U296 ( .A1(din[42]), .A2(n221), .B1(n222), .B2(n311), .C1(
        dout_eins[42]), .C2(n307), .O(din_eins[42]) );
  NR2 U297 ( .I1(din[42]), .I2(n91), .O(n222) );
  OAI12S U298 ( .B1(iv[42]), .B2(n339), .A1(n6), .O(n221) );
  AO222 U299 ( .A1(din[34]), .A2(n239), .B1(n240), .B2(n312), .C1(
        dout_eins[34]), .C2(n308), .O(din_eins[34]) );
  NR2 U300 ( .I1(din[34]), .I2(n109), .O(n240) );
  OAI12S U301 ( .B1(iv[34]), .B2(n337), .A1(n8), .O(n239) );
  AO222 U302 ( .A1(din[26]), .A2(n257), .B1(n258), .B2(n312), .C1(
        dout_eins[26]), .C2(n308), .O(din_eins[26]) );
  NR2 U303 ( .I1(din[26]), .I2(n127), .O(n258) );
  OAI12S U304 ( .B1(iv[26]), .B2(n336), .A1(n9), .O(n257) );
  AO222 U305 ( .A1(din[18]), .A2(n275), .B1(n276), .B2(n313), .C1(
        dout_eins[18]), .C2(n309), .O(din_eins[18]) );
  NR2 U306 ( .I1(din[18]), .I2(n145), .O(n276) );
  OAI12S U307 ( .B1(iv[18]), .B2(n335), .A1(n33), .O(n275) );
  AO222 U308 ( .A1(din[10]), .A2(n291), .B1(n292), .B2(n313), .C1(
        dout_eins[10]), .C2(n309), .O(din_eins[10]) );
  NR2 U309 ( .I1(din[10]), .I2(n161), .O(n292) );
  OAI12S U310 ( .B1(iv[10]), .B2(n334), .A1(n34), .O(n291) );
  AO222 U311 ( .A1(din[2]), .A2(n249), .B1(n250), .B2(n312), .C1(dout_eins[2]), 
        .C2(n308), .O(din_eins[2]) );
  NR2 U312 ( .I1(din[2]), .I2(n119), .O(n250) );
  OAI12S U313 ( .B1(iv[2]), .B2(n337), .A1(n8), .O(n249) );
  AO222 U314 ( .A1(din[60]), .A2(n181), .B1(n182), .B2(n310), .C1(
        dout_eins[60]), .C2(n306), .O(din_eins[60]) );
  NR2 U315 ( .I1(din[60]), .I2(n51), .O(n182) );
  OAI12S U316 ( .B1(iv[60]), .B2(n342), .A1(n3), .O(n181) );
  AO222 U317 ( .A1(din[52]), .A2(n199), .B1(n200), .B2(n311), .C1(
        dout_eins[52]), .C2(n307), .O(din_eins[52]) );
  NR2 U318 ( .I1(din[52]), .I2(n69), .O(n200) );
  OAI12S U319 ( .B1(iv[52]), .B2(n340), .A1(n4), .O(n199) );
  AO222 U320 ( .A1(din[44]), .A2(n217), .B1(n218), .B2(n311), .C1(
        dout_eins[44]), .C2(n307), .O(din_eins[44]) );
  NR2 U321 ( .I1(din[44]), .I2(n87), .O(n218) );
  OAI12S U322 ( .B1(iv[44]), .B2(n339), .A1(n6), .O(n217) );
  AO222 U323 ( .A1(din[36]), .A2(n235), .B1(n236), .B2(n312), .C1(
        dout_eins[36]), .C2(n308), .O(din_eins[36]) );
  NR2 U324 ( .I1(din[36]), .I2(n105), .O(n236) );
  OAI12S U325 ( .B1(iv[36]), .B2(n338), .A1(n7), .O(n235) );
  AO222 U326 ( .A1(din[28]), .A2(n253), .B1(n254), .B2(n312), .C1(
        dout_eins[28]), .C2(n308), .O(din_eins[28]) );
  NR2 U327 ( .I1(din[28]), .I2(n123), .O(n254) );
  OAI12S U328 ( .B1(iv[28]), .B2(n336), .A1(n9), .O(n253) );
  AO222 U329 ( .A1(din[20]), .A2(n269), .B1(n270), .B2(n313), .C1(
        dout_eins[20]), .C2(n309), .O(din_eins[20]) );
  NR2 U330 ( .I1(din[20]), .I2(n139), .O(n270) );
  OAI12S U331 ( .B1(iv[20]), .B2(n335), .A1(n26), .O(n269) );
  AO222 U332 ( .A1(din[12]), .A2(n287), .B1(n288), .B2(n313), .C1(
        dout_eins[12]), .C2(n309), .O(din_eins[12]) );
  NR2 U333 ( .I1(din[12]), .I2(n157), .O(n288) );
  OAI12S U334 ( .B1(iv[12]), .B2(n334), .A1(n34), .O(n287) );
  AO222 U335 ( .A1(din[4]), .A2(n205), .B1(n206), .B2(n311), .C1(dout_eins[4]), 
        .C2(n307), .O(din_eins[4]) );
  NR2 U336 ( .I1(din[4]), .I2(n75), .O(n206) );
  OAI12S U337 ( .B1(iv[4]), .B2(n340), .A1(n5), .O(n205) );
  AO222 U338 ( .A1(din[62]), .A2(n177), .B1(n178), .B2(n310), .C1(
        dout_eins[62]), .C2(n306), .O(din_eins[62]) );
  NR2 U339 ( .I1(din[62]), .I2(n47), .O(n178) );
  OAI12S U340 ( .B1(iv[62]), .B2(n342), .A1(n2), .O(n177) );
  AO222 U341 ( .A1(din[54]), .A2(n195), .B1(n196), .B2(n310), .C1(
        dout_eins[54]), .C2(n306), .O(din_eins[54]) );
  NR2 U342 ( .I1(din[54]), .I2(n65), .O(n196) );
  OAI12S U343 ( .B1(iv[54]), .B2(n341), .A1(n4), .O(n195) );
  AO222 U344 ( .A1(din[46]), .A2(n213), .B1(n214), .B2(n311), .C1(
        dout_eins[46]), .C2(n307), .O(din_eins[46]) );
  NR2 U345 ( .I1(din[46]), .I2(n83), .O(n214) );
  OAI12S U346 ( .B1(iv[46]), .B2(n339), .A1(n5), .O(n213) );
  AO222 U347 ( .A1(din[38]), .A2(n231), .B1(n232), .B2(n312), .C1(
        dout_eins[38]), .C2(n308), .O(din_eins[38]) );
  NR2 U348 ( .I1(din[38]), .I2(n101), .O(n232) );
  OAI12S U349 ( .B1(iv[38]), .B2(n338), .A1(n7), .O(n231) );
  AO222 U350 ( .A1(din[30]), .A2(n247), .B1(n248), .B2(n312), .C1(
        dout_eins[30]), .C2(n308), .O(din_eins[30]) );
  NR2 U351 ( .I1(din[30]), .I2(n117), .O(n248) );
  OAI12S U352 ( .B1(iv[30]), .B2(n337), .A1(n8), .O(n247) );
  AO222 U353 ( .A1(din[22]), .A2(n265), .B1(n266), .B2(n313), .C1(
        dout_eins[22]), .C2(n309), .O(din_eins[22]) );
  NR2 U354 ( .I1(din[22]), .I2(n135), .O(n266) );
  OAI12S U355 ( .B1(iv[22]), .B2(n335), .A1(n26), .O(n265) );
  AO222 U356 ( .A1(din[14]), .A2(n283), .B1(n284), .B2(n313), .C1(
        dout_eins[14]), .C2(n309), .O(din_eins[14]) );
  NR2 U357 ( .I1(din[14]), .I2(n153), .O(n284) );
  OAI12S U358 ( .B1(iv[14]), .B2(n334), .A1(n33), .O(n283) );
  AO222 U359 ( .A1(din[6]), .A2(n173), .B1(n174), .B2(n310), .C1(dout_eins[6]), 
        .C2(n306), .O(din_eins[6]) );
  NR2 U360 ( .I1(din[6]), .I2(n43), .O(n174) );
  OAI12S U361 ( .B1(iv[6]), .B2(n342), .A1(n2), .O(n173) );
  XNR2 U362 ( .I1(n301), .I2(round[1]), .O(n23) );
  OAI12S U363 ( .B1(n302), .B2(n303), .A1(n300), .O(n301) );
  OAI112S U364 ( .C1(n343), .C2(n11), .A1(n12), .B1(n13), .O(n304) );
  INV2 U365 ( .I(dt_sel), .O(n11) );
  ND2 U366 ( .I1(test_so), .I2(n14), .O(n13) );
  OAI112S U367 ( .C1(n15), .C2(n16), .A1(n17), .B1(n12), .O(n305) );
  ND3 U368 ( .I1(dt_sel), .I2(n16), .I3(n15), .O(n17) );
  INV2 U369 ( .I(n14), .O(n15) );
  INV2 U370 ( .I(edr[0]), .O(n302) );
  XOR2 U371 ( .I1(dout_eins[46]), .I2(n82), .O(dout[46]) );
  NR2 U372 ( .I1(n316), .I2(n83), .O(n82) );
  XOR2 U373 ( .I1(dout_eins[47]), .I2(n80), .O(dout[47]) );
  NR2 U374 ( .I1(n316), .I2(n81), .O(n80) );
  XOR2 U375 ( .I1(dout_eins[48]), .I2(n78), .O(dout[48]) );
  NR2 U376 ( .I1(n316), .I2(n79), .O(n78) );
  XOR2 U377 ( .I1(dout_eins[49]), .I2(n76), .O(dout[49]) );
  NR2 U378 ( .I1(n316), .I2(n77), .O(n76) );
  XOR2 U379 ( .I1(dout_eins[50]), .I2(n72), .O(dout[50]) );
  NR2 U380 ( .I1(n316), .I2(n73), .O(n72) );
  XOR2 U381 ( .I1(dout_eins[51]), .I2(n70), .O(dout[51]) );
  NR2 U382 ( .I1(n316), .I2(n71), .O(n70) );
  XOR2 U383 ( .I1(dout_eins[1]), .I2(n140), .O(dout[1]) );
  NR2 U384 ( .I1(n320), .I2(n141), .O(n140) );
  XOR2 U385 ( .I1(dout_eins[32]), .I2(n112), .O(dout[32]) );
  NR2 U386 ( .I1(n318), .I2(n113), .O(n112) );
  XOR2 U387 ( .I1(dout_eins[33]), .I2(n110), .O(dout[33]) );
  NR2 U388 ( .I1(n318), .I2(n111), .O(n110) );
  XOR2 U389 ( .I1(dout_eins[34]), .I2(n108), .O(dout[34]) );
  NR2 U390 ( .I1(n318), .I2(n109), .O(n108) );
  XOR2 U391 ( .I1(dout_eins[35]), .I2(n106), .O(dout[35]) );
  NR2 U392 ( .I1(n318), .I2(n107), .O(n106) );
  XOR2 U393 ( .I1(dout_eins[36]), .I2(n104), .O(dout[36]) );
  NR2 U394 ( .I1(n318), .I2(n105), .O(n104) );
  XOR2 U395 ( .I1(dout_eins[37]), .I2(n102), .O(dout[37]) );
  NR2 U396 ( .I1(n318), .I2(n103), .O(n102) );
  XOR2 U397 ( .I1(dout_eins[38]), .I2(n100), .O(dout[38]) );
  NR2 U398 ( .I1(n318), .I2(n101), .O(n100) );
  XOR2 U399 ( .I1(dout_eins[39]), .I2(n98), .O(dout[39]) );
  NR2 U400 ( .I1(n317), .I2(n99), .O(n98) );
  XOR2 U401 ( .I1(dout_eins[40]), .I2(n94), .O(dout[40]) );
  NR2 U402 ( .I1(n317), .I2(n95), .O(n94) );
  XOR2 U403 ( .I1(dout_eins[41]), .I2(n92), .O(dout[41]) );
  NR2 U404 ( .I1(n317), .I2(n93), .O(n92) );
  XOR2 U405 ( .I1(dout_eins[42]), .I2(n90), .O(dout[42]) );
  NR2 U406 ( .I1(n317), .I2(n91), .O(n90) );
  XOR2 U407 ( .I1(dout_eins[52]), .I2(n68), .O(dout[52]) );
  NR2 U408 ( .I1(n316), .I2(n69), .O(n68) );
  XOR2 U409 ( .I1(dout_eins[53]), .I2(n66), .O(dout[53]) );
  NR2 U410 ( .I1(n315), .I2(n67), .O(n66) );
  XOR2 U411 ( .I1(dout_eins[54]), .I2(n64), .O(dout[54]) );
  NR2 U412 ( .I1(n315), .I2(n65), .O(n64) );
  XOR2 U413 ( .I1(dout_eins[55]), .I2(n62), .O(dout[55]) );
  NR2 U414 ( .I1(n315), .I2(n63), .O(n62) );
  XOR2 U415 ( .I1(dout_eins[56]), .I2(n60), .O(dout[56]) );
  NR2 U416 ( .I1(n315), .I2(n61), .O(n60) );
  XOR2 U417 ( .I1(dout_eins[57]), .I2(n58), .O(dout[57]) );
  NR2 U418 ( .I1(n315), .I2(n59), .O(n58) );
  XOR2 U419 ( .I1(dout_eins[58]), .I2(n56), .O(dout[58]) );
  NR2 U420 ( .I1(n315), .I2(n57), .O(n56) );
  XOR2 U421 ( .I1(dout_eins[59]), .I2(n54), .O(dout[59]) );
  NR2 U422 ( .I1(n315), .I2(n55), .O(n54) );
  XOR2 U423 ( .I1(dout_eins[60]), .I2(n50), .O(dout[60]) );
  NR2 U424 ( .I1(n314), .I2(n51), .O(n50) );
  XOR2 U425 ( .I1(dout_eins[61]), .I2(n48), .O(dout[61]) );
  NR2 U426 ( .I1(n314), .I2(n49), .O(n48) );
  XOR2 U427 ( .I1(dout_eins[62]), .I2(n46), .O(dout[62]) );
  NR2 U428 ( .I1(n314), .I2(n47), .O(n46) );
  XOR2 U429 ( .I1(dout_eins[63]), .I2(n44), .O(dout[63]) );
  NR2 U430 ( .I1(n314), .I2(n45), .O(n44) );
  XOR2 U431 ( .I1(dout_eins[0]), .I2(n162), .O(dout[0]) );
  NR2 U432 ( .I1(n321), .I2(n163), .O(n162) );
  XOR2 U433 ( .I1(dout_eins[2]), .I2(n118), .O(dout[2]) );
  NR2 U434 ( .I1(n319), .I2(n119), .O(n118) );
  XOR2 U435 ( .I1(dout_eins[3]), .I2(n96), .O(dout[3]) );
  NR2 U436 ( .I1(n317), .I2(n97), .O(n96) );
  XOR2 U437 ( .I1(dout_eins[4]), .I2(n74), .O(dout[4]) );
  NR2 U438 ( .I1(n316), .I2(n75), .O(n74) );
  XOR2 U439 ( .I1(dout_eins[5]), .I2(n52), .O(dout[5]) );
  NR2 U440 ( .I1(n315), .I2(n53), .O(n52) );
  XOR2 U441 ( .I1(dout_eins[6]), .I2(n42), .O(dout[6]) );
  NR2 U442 ( .I1(n314), .I2(n43), .O(n42) );
  XOR2 U443 ( .I1(dout_eins[7]), .I2(n40), .O(dout[7]) );
  NR2 U444 ( .I1(n314), .I2(n41), .O(n40) );
  XOR2 U445 ( .I1(dout_eins[8]), .I2(n38), .O(dout[8]) );
  NR2 U446 ( .I1(n314), .I2(n39), .O(n38) );
  XOR2 U447 ( .I1(dout_eins[9]), .I2(n35), .O(dout[9]) );
  NR2 U448 ( .I1(n314), .I2(n37), .O(n35) );
  XOR2 U449 ( .I1(dout_eins[10]), .I2(n160), .O(dout[10]) );
  NR2 U450 ( .I1(n321), .I2(n161), .O(n160) );
  XOR2 U451 ( .I1(dout_eins[11]), .I2(n158), .O(dout[11]) );
  NR2 U452 ( .I1(n321), .I2(n159), .O(n158) );
  XOR2 U453 ( .I1(dout_eins[12]), .I2(n156), .O(dout[12]) );
  NR2 U454 ( .I1(n321), .I2(n157), .O(n156) );
  XOR2 U455 ( .I1(dout_eins[13]), .I2(n154), .O(dout[13]) );
  NR2 U456 ( .I1(n321), .I2(n155), .O(n154) );
  XOR2 U457 ( .I1(dout_eins[14]), .I2(n152), .O(dout[14]) );
  NR2 U458 ( .I1(n321), .I2(n153), .O(n152) );
  XOR2 U459 ( .I1(dout_eins[15]), .I2(n150), .O(dout[15]) );
  NR2 U460 ( .I1(n321), .I2(n151), .O(n150) );
  XOR2 U461 ( .I1(dout_eins[16]), .I2(n148), .O(dout[16]) );
  NR2 U462 ( .I1(n321), .I2(n149), .O(n148) );
  XOR2 U463 ( .I1(dout_eins[17]), .I2(n146), .O(dout[17]) );
  NR2 U464 ( .I1(n320), .I2(n147), .O(n146) );
  XOR2 U465 ( .I1(dout_eins[18]), .I2(n144), .O(dout[18]) );
  NR2 U466 ( .I1(n320), .I2(n145), .O(n144) );
  XOR2 U467 ( .I1(dout_eins[19]), .I2(n142), .O(dout[19]) );
  NR2 U468 ( .I1(n320), .I2(n143), .O(n142) );
  XOR2 U469 ( .I1(dout_eins[20]), .I2(n138), .O(dout[20]) );
  NR2 U470 ( .I1(n320), .I2(n139), .O(n138) );
  XOR2 U471 ( .I1(dout_eins[21]), .I2(n136), .O(dout[21]) );
  NR2 U472 ( .I1(n320), .I2(n137), .O(n136) );
  XOR2 U473 ( .I1(dout_eins[22]), .I2(n134), .O(dout[22]) );
  NR2 U474 ( .I1(n320), .I2(n135), .O(n134) );
  XOR2 U475 ( .I1(dout_eins[23]), .I2(n132), .O(dout[23]) );
  NR2 U476 ( .I1(n320), .I2(n133), .O(n132) );
  XOR2 U477 ( .I1(dout_eins[24]), .I2(n130), .O(dout[24]) );
  NR2 U478 ( .I1(n319), .I2(n131), .O(n130) );
  XOR2 U479 ( .I1(dout_eins[25]), .I2(n128), .O(dout[25]) );
  NR2 U480 ( .I1(n319), .I2(n129), .O(n128) );
  XOR2 U481 ( .I1(dout_eins[26]), .I2(n126), .O(dout[26]) );
  NR2 U482 ( .I1(n319), .I2(n127), .O(n126) );
  XOR2 U483 ( .I1(dout_eins[27]), .I2(n124), .O(dout[27]) );
  NR2 U484 ( .I1(n319), .I2(n125), .O(n124) );
  XOR2 U485 ( .I1(dout_eins[28]), .I2(n122), .O(dout[28]) );
  NR2 U486 ( .I1(n319), .I2(n123), .O(n122) );
  XOR2 U487 ( .I1(dout_eins[29]), .I2(n120), .O(dout[29]) );
  NR2 U488 ( .I1(n319), .I2(n121), .O(n120) );
  XOR2 U489 ( .I1(dout_eins[30]), .I2(n116), .O(dout[30]) );
  NR2 U490 ( .I1(n319), .I2(n117), .O(n116) );
  XOR2 U491 ( .I1(dout_eins[31]), .I2(n114), .O(dout[31]) );
  NR2 U492 ( .I1(n318), .I2(n115), .O(n114) );
  INV2 U493 ( .I(edr[1]), .O(n303) );
  XOR2 U494 ( .I1(dout_eins[43]), .I2(n88), .O(dout[43]) );
  NR2 U495 ( .I1(n317), .I2(n89), .O(n88) );
  XOR2 U496 ( .I1(dout_eins[44]), .I2(n86), .O(dout[44]) );
  NR2 U497 ( .I1(n317), .I2(n87), .O(n86) );
  XOR2 U498 ( .I1(dout_eins[45]), .I2(n84), .O(dout[45]) );
  NR2 U499 ( .I1(n317), .I2(n85), .O(n84) );
  XNR2 U500 ( .I1(encrypt_whole), .I2(n1), .O(encrypt_eins) );
  ND3T U501 ( .I1(iv_sel), .I2(encrypt_whole), .I3(mode_sel), .O(n36) );
  XOR2 U502 ( .I1(n300), .I2(round[2]), .O(n18) );
  XOR2 U503 ( .I1(n300), .I2(round[3]), .O(n19) );
  XOR2 U504 ( .I1(edr[0]), .I2(round[0]), .O(n21) );
  OAI12S U505 ( .B1(n298), .B2(n299), .A1(n12), .O(N31) );
  ND3 U506 ( .I1(n19), .I2(dt_sel), .I3(n18), .O(n299) );
  ND3 U507 ( .I1(n21), .I2(n23), .I3(test_so), .O(n298) );
  INV2 U508 ( .I(iv[56]), .O(n61) );
  INV2 U509 ( .I(iv[48]), .O(n79) );
  INV2 U510 ( .I(iv[40]), .O(n95) );
  INV2 U511 ( .I(iv[32]), .O(n113) );
  INV2 U512 ( .I(iv[24]), .O(n131) );
  INV2 U513 ( .I(iv[16]), .O(n149) );
  INV2 U514 ( .I(iv[8]), .O(n39) );
  INV2 U515 ( .I(iv[0]), .O(n163) );
  INV2 U516 ( .I(iv[58]), .O(n57) );
  INV2 U517 ( .I(iv[50]), .O(n73) );
  INV2 U518 ( .I(iv[42]), .O(n91) );
  INV2 U519 ( .I(iv[34]), .O(n109) );
  INV2 U520 ( .I(iv[26]), .O(n127) );
  INV2 U521 ( .I(iv[18]), .O(n145) );
  INV2 U522 ( .I(iv[10]), .O(n161) );
  INV2 U523 ( .I(iv[2]), .O(n119) );
  INV2 U524 ( .I(iv[60]), .O(n51) );
  INV2 U525 ( .I(iv[52]), .O(n69) );
  INV2 U526 ( .I(iv[44]), .O(n87) );
  INV2 U527 ( .I(iv[36]), .O(n105) );
  INV2 U528 ( .I(iv[28]), .O(n123) );
  INV2 U529 ( .I(iv[20]), .O(n139) );
  INV2 U530 ( .I(iv[12]), .O(n157) );
  INV2 U531 ( .I(iv[4]), .O(n75) );
  INV2 U532 ( .I(iv[62]), .O(n47) );
  INV2 U533 ( .I(iv[54]), .O(n65) );
  INV2 U534 ( .I(iv[46]), .O(n83) );
  INV2 U535 ( .I(iv[38]), .O(n101) );
  INV2 U536 ( .I(iv[30]), .O(n117) );
  INV2 U537 ( .I(iv[22]), .O(n135) );
  INV2 U538 ( .I(iv[14]), .O(n153) );
  INV2 U539 ( .I(iv[6]), .O(n43) );
  INV2 U540 ( .I(din_valid_whole), .O(n12) );
  QDFZRBS din_valid_eins_reg ( .D(N31), .TD(dout_eins[7]), .SEL(test_se), .CK(
        hclk), .RB(hresetn), .Q(din_valid_eins) );
  QDFZRBS flag_reg_1 ( .D(n304), .TD(flag_0_), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(test_so) );
  QDFZRBS flag_reg_0 ( .D(n305), .TD(din_valid_eins), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(flag_0_) );
endmodule


module des_dat ( POR, hresetn, clrptr, hclk, rd, wr, deswr, data, data_all, 
        full_pulse, q, q_all, test_mode, test_se, test_si, test_so );
  input [31:0] data;
  input [63:0] data_all;
  output [31:0] q;
  output [63:0] q_all;
  input POR, hresetn, clrptr, hclk, rd, wr, deswr, test_mode, test_se, test_si;
  output full_pulse, test_so;
  wire   N4, N9, N11, N13, N15, N17, N19, N21, N23, N25, N27, N29, N31, N33,
         N35, N37, N39, N41, N43, N45, N47, N49, N51, N53, N55, N57, N59, N61,
         N63, N65, N67, N69, N70, N71, N73, N75, N77, N79, N81, N83, N85, N87,
         N89, N91, N93, N95, N97, N99, N101, N103, N105, N107, N109, N111,
         N113, N115, N117, N119, N121, N123, N125, N127, N129, N131, N133,
         N134, N135, full, N161, full_delay, N162, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195,
         CLKGATING_hclk_POWERGATING_hclk_N134_0_0, net1811,
         CLKGATING_hclk_POWERGATING_hclk_N70_0_0, net1816, n6, n7, n8, n9, n10,
         n11, n12, n13, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n1, n2, n3, n4, n5, n14, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n78;
  wire   [1:0] ptr;

  POWERMODULE_HIGH_des_dat_0_1 POWERGATING_hclk_N134_0 ( .CLK(hclk), .EN(N134), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .TE(n70), .ENOBS(
        net1811) );
  POWERMODULE_HIGH_des_dat_0_0 POWERGATING_hclk_N70_0 ( .CLK(hclk), .EN(N70), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .TE(n70), .ENOBS(
        net1816) );
  SNPS_CLOCK_GATE_OBS_des_dat clk_gate_obs ( .TE(n70), .net1811(net1811), 
        .net1816(net1816), .hclk(hclk), .test_se(test_se), .test_si(test_si), 
        .test_so(n78) );
  BUF1 U3 ( .I(test_mode), .O(n70) );
  INV3 U4 ( .I(n74), .O(n71) );
  INV3 U5 ( .I(n75), .O(n72) );
  INV2 U6 ( .I(n74), .O(n73) );
  BUF1 U7 ( .I(n21), .O(n61) );
  BUF2 U8 ( .I(n21), .O(n60) );
  BUF2 U9 ( .I(n21), .O(n3) );
  BUF2 U10 ( .I(n21), .O(n4) );
  BUF2 U11 ( .I(n21), .O(n5) );
  BUF2 U12 ( .I(n21), .O(n14) );
  BUF2 U13 ( .I(n21), .O(n59) );
  BUF1 U14 ( .I(n76), .O(n74) );
  BUF1 U15 ( .I(n76), .O(n75) );
  BUF2 U16 ( .I(n12), .O(n62) );
  INV2 U17 ( .I(n36), .O(n21) );
  BUF2 U18 ( .I(n12), .O(n68) );
  BUF2 U19 ( .I(n12), .O(n63) );
  BUF2 U20 ( .I(n12), .O(n64) );
  BUF2 U21 ( .I(n12), .O(n65) );
  BUF2 U22 ( .I(n12), .O(n66) );
  BUF2 U23 ( .I(n12), .O(n67) );
  BUF1 U24 ( .I(n12), .O(n69) );
  INV2 U25 ( .I(rd), .O(n76) );
  INV2 U26 ( .I(wr), .O(n12) );
  ND2 U27 ( .I1(deswr), .I2(n62), .O(n36) );
  INV2 U28 ( .I(clrptr), .O(n7) );
  ND2 U29 ( .I1(wr), .I2(n11), .O(n8) );
  AN2 U30 ( .I1(N195), .I2(n71), .O(q[0]) );
  MUX2 U31 ( .A(q_all[0]), .B(q_all[32]), .S(n1), .O(N195) );
  AN2 U32 ( .I1(N194), .I2(n71), .O(q[1]) );
  MUX2 U33 ( .A(q_all[1]), .B(q_all[33]), .S(n1), .O(N194) );
  AN2 U34 ( .I1(N193), .I2(n72), .O(q[2]) );
  MUX2 U35 ( .A(q_all[2]), .B(q_all[34]), .S(n1), .O(N193) );
  AN2 U36 ( .I1(N192), .I2(n72), .O(q[3]) );
  MUX2 U37 ( .A(q_all[3]), .B(q_all[35]), .S(n1), .O(N192) );
  AN2 U38 ( .I1(N191), .I2(n72), .O(q[4]) );
  MUX2 U39 ( .A(q_all[4]), .B(q_all[36]), .S(n1), .O(N191) );
  AN2 U40 ( .I1(N190), .I2(n72), .O(q[5]) );
  MUX2 U41 ( .A(q_all[5]), .B(q_all[37]), .S(n1), .O(N190) );
  AN2 U42 ( .I1(N189), .I2(n72), .O(q[6]) );
  MUX2 U43 ( .A(q_all[6]), .B(q_all[38]), .S(n1), .O(N189) );
  AN2 U44 ( .I1(N188), .I2(n72), .O(q[7]) );
  MUX2 U45 ( .A(q_all[7]), .B(q_all[39]), .S(n1), .O(N188) );
  AN2 U46 ( .I1(N185), .I2(n71), .O(q[10]) );
  MUX2 U47 ( .A(q_all[10]), .B(q_all[42]), .S(n1), .O(N185) );
  AN2 U48 ( .I1(N184), .I2(n71), .O(q[11]) );
  MUX2 U49 ( .A(q_all[11]), .B(q_all[43]), .S(n1), .O(N184) );
  AN2 U50 ( .I1(N183), .I2(n71), .O(q[12]) );
  MUX2 U51 ( .A(q_all[12]), .B(q_all[44]), .S(n1), .O(N183) );
  AN2 U52 ( .I1(N182), .I2(n71), .O(q[13]) );
  MUX2 U53 ( .A(q_all[13]), .B(q_all[45]), .S(n1), .O(N182) );
  AN2 U54 ( .I1(N181), .I2(n71), .O(q[14]) );
  MUX2 U55 ( .A(q_all[14]), .B(q_all[46]), .S(n1), .O(N181) );
  AN2 U56 ( .I1(N180), .I2(n72), .O(q[15]) );
  MUX2 U57 ( .A(q_all[15]), .B(q_all[47]), .S(n1), .O(N180) );
  AN2 U58 ( .I1(N179), .I2(n71), .O(q[16]) );
  MUX2 U59 ( .A(q_all[16]), .B(q_all[48]), .S(n2), .O(N179) );
  AN2 U60 ( .I1(N178), .I2(n71), .O(q[17]) );
  MUX2 U61 ( .A(q_all[17]), .B(q_all[49]), .S(n2), .O(N178) );
  AN2 U62 ( .I1(N177), .I2(n71), .O(q[18]) );
  MUX2 U63 ( .A(q_all[18]), .B(q_all[50]), .S(n2), .O(N177) );
  AN2 U64 ( .I1(N176), .I2(n71), .O(q[19]) );
  MUX2 U65 ( .A(q_all[19]), .B(q_all[51]), .S(n2), .O(N176) );
  AN2 U66 ( .I1(N175), .I2(n71), .O(q[20]) );
  MUX2 U67 ( .A(q_all[20]), .B(q_all[52]), .S(n2), .O(N175) );
  AN2 U68 ( .I1(N174), .I2(n71), .O(q[21]) );
  MUX2 U69 ( .A(q_all[21]), .B(q_all[53]), .S(n2), .O(N174) );
  AN2 U70 ( .I1(N173), .I2(n71), .O(q[22]) );
  MUX2 U71 ( .A(q_all[22]), .B(q_all[54]), .S(n2), .O(N173) );
  AN2 U72 ( .I1(N172), .I2(n72), .O(q[23]) );
  MUX2 U73 ( .A(q_all[23]), .B(q_all[55]), .S(n2), .O(N172) );
  AN2 U74 ( .I1(N171), .I2(n72), .O(q[24]) );
  MUX2 U75 ( .A(q_all[24]), .B(q_all[56]), .S(n2), .O(N171) );
  AN2 U76 ( .I1(N170), .I2(n72), .O(q[25]) );
  MUX2 U77 ( .A(q_all[25]), .B(q_all[57]), .S(n2), .O(N170) );
  AN2 U78 ( .I1(N169), .I2(n72), .O(q[26]) );
  MUX2 U79 ( .A(q_all[26]), .B(q_all[58]), .S(n2), .O(N169) );
  AN2 U80 ( .I1(N168), .I2(n72), .O(q[27]) );
  MUX2 U81 ( .A(q_all[27]), .B(q_all[59]), .S(n2), .O(N168) );
  AN2 U82 ( .I1(N167), .I2(n72), .O(q[28]) );
  MUX2 U83 ( .A(q_all[28]), .B(q_all[60]), .S(n2), .O(N167) );
  AN2 U84 ( .I1(N166), .I2(n72), .O(q[29]) );
  MUX2 U85 ( .A(q_all[29]), .B(q_all[61]), .S(n2), .O(N166) );
  AN2 U86 ( .I1(N165), .I2(n72), .O(q[30]) );
  MUX2 U87 ( .A(q_all[30]), .B(q_all[62]), .S(n2), .O(N165) );
  AN2 U88 ( .I1(N164), .I2(n72), .O(q[31]) );
  MUX2 U89 ( .A(q_all[31]), .B(q_all[63]), .S(n2), .O(N164) );
  AN2 U90 ( .I1(N187), .I2(n73), .O(q[8]) );
  MUX2 U91 ( .A(q_all[8]), .B(q_all[40]), .S(n1), .O(N187) );
  AN2 U92 ( .I1(n73), .I2(N186), .O(q[9]) );
  MUX2 U93 ( .A(q_all[9]), .B(q_all[41]), .S(n1), .O(N186) );
  BUF2 U94 ( .I(N4), .O(n1) );
  BUF2 U95 ( .I(N4), .O(n2) );
  AO12 U96 ( .B1(wr), .B2(test_so), .A1(n61), .O(N134) );
  OAI12S U97 ( .B1(test_so), .B2(n62), .A1(n36), .O(N70) );
  MOAI1 U98 ( .A1(n62), .A2(n53), .B1(data_all[46]), .B2(n14), .O(N101) );
  MOAI1 U99 ( .A1(n62), .A2(n52), .B1(data_all[47]), .B2(n3), .O(N103) );
  MOAI1 U100 ( .A1(n62), .A2(n51), .B1(data_all[48]), .B2(n3), .O(N105) );
  MOAI1 U101 ( .A1(n62), .A2(n50), .B1(data_all[49]), .B2(n3), .O(N107) );
  MOAI1 U102 ( .A1(n62), .A2(n49), .B1(data_all[50]), .B2(n3), .O(N109) );
  MOAI1 U103 ( .A1(n62), .A2(n48), .B1(data_all[51]), .B2(n3), .O(N111) );
  MOAI1 U104 ( .A1(n62), .A2(n34), .B1(data_all[1]), .B2(n3), .O(N11) );
  MOAI1 U105 ( .A1(n67), .A2(n26), .B1(data_all[32]), .B2(n60), .O(N73) );
  MOAI1 U106 ( .A1(n67), .A2(n34), .B1(data_all[33]), .B2(n60), .O(N75) );
  MOAI1 U107 ( .A1(n67), .A2(n33), .B1(data_all[34]), .B2(n60), .O(N77) );
  MOAI1 U108 ( .A1(n68), .A2(n32), .B1(data_all[35]), .B2(n60), .O(N79) );
  MOAI1 U109 ( .A1(n68), .A2(n31), .B1(data_all[36]), .B2(n60), .O(N81) );
  MOAI1 U110 ( .A1(n68), .A2(n30), .B1(data_all[37]), .B2(n60), .O(N83) );
  MOAI1 U111 ( .A1(n68), .A2(n29), .B1(data_all[38]), .B2(n60), .O(N85) );
  MOAI1 U112 ( .A1(n68), .A2(n28), .B1(data_all[39]), .B2(n60), .O(N87) );
  MOAI1 U113 ( .A1(n68), .A2(n27), .B1(data_all[40]), .B2(n60), .O(N89) );
  MOAI1 U114 ( .A1(n68), .A2(n25), .B1(data_all[41]), .B2(n61), .O(N91) );
  MOAI1 U115 ( .A1(n68), .A2(n24), .B1(data_all[42]), .B2(n61), .O(N93) );
  MOAI1 U116 ( .A1(n63), .A2(n47), .B1(data_all[52]), .B2(n3), .O(N113) );
  MOAI1 U117 ( .A1(n63), .A2(n46), .B1(data_all[53]), .B2(n3), .O(N115) );
  MOAI1 U118 ( .A1(n63), .A2(n45), .B1(data_all[54]), .B2(n3), .O(N117) );
  MOAI1 U119 ( .A1(n63), .A2(n44), .B1(data_all[55]), .B2(n4), .O(N119) );
  MOAI1 U120 ( .A1(n63), .A2(n43), .B1(data_all[56]), .B2(n4), .O(N121) );
  MOAI1 U121 ( .A1(n63), .A2(n42), .B1(data_all[57]), .B2(n4), .O(N123) );
  MOAI1 U122 ( .A1(n63), .A2(n41), .B1(data_all[58]), .B2(n4), .O(N125) );
  MOAI1 U123 ( .A1(n63), .A2(n40), .B1(data_all[59]), .B2(n4), .O(N127) );
  MOAI1 U124 ( .A1(n65), .A2(n39), .B1(data_all[60]), .B2(n4), .O(N129) );
  MOAI1 U125 ( .A1(n64), .A2(n38), .B1(data_all[61]), .B2(n4), .O(N131) );
  MOAI1 U126 ( .A1(n64), .A2(n37), .B1(data_all[62]), .B2(n4), .O(N133) );
  MOAI1 U127 ( .A1(n64), .A2(n35), .B1(data_all[63]), .B2(n4), .O(N135) );
  MOAI1 U128 ( .A1(n68), .A2(n26), .B1(data_all[0]), .B2(n60), .O(N9) );
  MOAI1 U129 ( .A1(n63), .A2(n33), .B1(data_all[2]), .B2(n4), .O(N13) );
  MOAI1 U130 ( .A1(n64), .A2(n32), .B1(data_all[3]), .B2(n5), .O(N15) );
  MOAI1 U131 ( .A1(n64), .A2(n31), .B1(data_all[4]), .B2(n5), .O(N17) );
  MOAI1 U132 ( .A1(n64), .A2(n30), .B1(data_all[5]), .B2(n5), .O(N19) );
  MOAI1 U133 ( .A1(n64), .A2(n29), .B1(data_all[6]), .B2(n5), .O(N21) );
  MOAI1 U134 ( .A1(n64), .A2(n28), .B1(data_all[7]), .B2(n5), .O(N23) );
  MOAI1 U135 ( .A1(n64), .A2(n27), .B1(data_all[8]), .B2(n5), .O(N25) );
  MOAI1 U136 ( .A1(n65), .A2(n25), .B1(data_all[9]), .B2(n5), .O(N27) );
  MOAI1 U137 ( .A1(n65), .A2(n24), .B1(data_all[10]), .B2(n5), .O(N29) );
  MOAI1 U138 ( .A1(n65), .A2(n23), .B1(data_all[11]), .B2(n5), .O(N31) );
  MOAI1 U139 ( .A1(n65), .A2(n22), .B1(data_all[12]), .B2(n5), .O(N33) );
  MOAI1 U140 ( .A1(n65), .A2(n20), .B1(data_all[13]), .B2(n14), .O(N35) );
  MOAI1 U141 ( .A1(n65), .A2(n53), .B1(data_all[14]), .B2(n14), .O(N37) );
  MOAI1 U142 ( .A1(n65), .A2(n52), .B1(data_all[15]), .B2(n14), .O(N39) );
  MOAI1 U143 ( .A1(n65), .A2(n51), .B1(data_all[16]), .B2(n14), .O(N41) );
  MOAI1 U144 ( .A1(n66), .A2(n50), .B1(data_all[17]), .B2(n14), .O(N43) );
  MOAI1 U145 ( .A1(n66), .A2(n49), .B1(data_all[18]), .B2(n14), .O(N45) );
  MOAI1 U146 ( .A1(n66), .A2(n48), .B1(data_all[19]), .B2(n14), .O(N47) );
  MOAI1 U147 ( .A1(n66), .A2(n47), .B1(data_all[20]), .B2(n14), .O(N49) );
  MOAI1 U148 ( .A1(n66), .A2(n46), .B1(data_all[21]), .B2(n14), .O(N51) );
  MOAI1 U149 ( .A1(n66), .A2(n45), .B1(data_all[22]), .B2(n59), .O(N53) );
  MOAI1 U150 ( .A1(n66), .A2(n44), .B1(data_all[23]), .B2(n59), .O(N55) );
  MOAI1 U151 ( .A1(n66), .A2(n43), .B1(data_all[24]), .B2(n59), .O(N57) );
  MOAI1 U152 ( .A1(n66), .A2(n42), .B1(data_all[25]), .B2(n59), .O(N59) );
  MOAI1 U153 ( .A1(n67), .A2(n41), .B1(data_all[26]), .B2(n59), .O(N61) );
  MOAI1 U154 ( .A1(n67), .A2(n40), .B1(data_all[27]), .B2(n59), .O(N63) );
  MOAI1 U155 ( .A1(n67), .A2(n39), .B1(data_all[28]), .B2(n59), .O(N65) );
  MOAI1 U156 ( .A1(n67), .A2(n38), .B1(data_all[29]), .B2(n59), .O(N67) );
  MOAI1 U157 ( .A1(n67), .A2(n37), .B1(data_all[30]), .B2(n59), .O(N69) );
  MOAI1 U158 ( .A1(n67), .A2(n35), .B1(data_all[31]), .B2(n59), .O(N71) );
  MOAI1 U159 ( .A1(n69), .A2(n23), .B1(data_all[43]), .B2(n61), .O(N95) );
  MOAI1 U160 ( .A1(n69), .A2(n22), .B1(data_all[44]), .B2(n61), .O(N97) );
  MOAI1 U161 ( .A1(n69), .A2(n20), .B1(data_all[45]), .B2(n3), .O(N99) );
  NR3P U162 ( .I1(n7), .I2(ptr[0]), .I3(n11), .O(N161) );
  NR2 U163 ( .I1(n15), .I2(n7), .O(n57) );
  XOR2 U164 ( .I1(n16), .I2(N4), .O(n15) );
  OAI12S U165 ( .B1(n17), .B2(ptr[1]), .A1(n71), .O(n16) );
  NR2 U166 ( .I1(wr), .I2(n13), .O(n17) );
  MOAI1 U167 ( .A1(n18), .A2(n7), .B1(N161), .B2(n71), .O(n58) );
  AOI13HS U168 ( .B1(n8), .B2(n75), .B3(ptr[0]), .A1(n19), .O(n18) );
  NR2 U169 ( .I1(ptr[0]), .I2(n8), .O(n19) );
  NR2 U170 ( .I1(n9), .I2(n7), .O(n56) );
  OA22 U171 ( .A1(n10), .A2(n11), .B1(n69), .B2(n13), .O(n9) );
  NR2 U172 ( .I1(ptr[0]), .I2(n74), .O(n10) );
  INV2 U173 ( .I(ptr[1]), .O(n11) );
  INV2 U174 ( .I(data[1]), .O(n34) );
  INV2 U175 ( .I(data[2]), .O(n33) );
  INV2 U176 ( .I(data[3]), .O(n32) );
  INV2 U177 ( .I(data[4]), .O(n31) );
  INV2 U178 ( .I(data[5]), .O(n30) );
  INV2 U179 ( .I(data[6]), .O(n29) );
  INV2 U180 ( .I(data[7]), .O(n28) );
  INV2 U181 ( .I(data[9]), .O(n25) );
  INV2 U182 ( .I(data[10]), .O(n24) );
  INV2 U183 ( .I(data[11]), .O(n23) );
  INV2 U184 ( .I(data[12]), .O(n22) );
  INV2 U185 ( .I(data[13]), .O(n20) );
  INV2 U186 ( .I(data[14]), .O(n53) );
  INV2 U187 ( .I(data[15]), .O(n52) );
  INV2 U188 ( .I(data[17]), .O(n50) );
  INV2 U189 ( .I(data[18]), .O(n49) );
  INV2 U190 ( .I(data[19]), .O(n48) );
  INV2 U191 ( .I(data[20]), .O(n47) );
  INV2 U192 ( .I(data[21]), .O(n46) );
  INV2 U193 ( .I(data[22]), .O(n45) );
  INV2 U194 ( .I(data[23]), .O(n44) );
  INV2 U195 ( .I(data[25]), .O(n42) );
  INV2 U196 ( .I(data[26]), .O(n41) );
  INV2 U197 ( .I(data[27]), .O(n40) );
  INV2 U198 ( .I(data[28]), .O(n39) );
  INV2 U199 ( .I(data[29]), .O(n38) );
  INV2 U200 ( .I(data[30]), .O(n37) );
  INV2 U201 ( .I(data[31]), .O(n35) );
  NR2 U202 ( .I1(n6), .I2(n7), .O(n55) );
  XOR2 U203 ( .I1(n8), .I2(test_so), .O(n6) );
  INV2 U204 ( .I(data[0]), .O(n26) );
  INV2 U205 ( .I(data[8]), .O(n27) );
  INV2 U206 ( .I(data[16]), .O(n51) );
  INV2 U207 ( .I(data[24]), .O(n43) );
  INV2 U208 ( .I(ptr[0]), .O(n13) );
  NR2 U209 ( .I1(full_delay), .I2(n54), .O(N162) );
  INV2 U210 ( .I(full), .O(n54) );
  QDFZRBS full_delay_reg ( .D(full), .TD(q_all[63]), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(full_delay) );
  QDFZRBS full_reg ( .D(N161), .TD(full_pulse), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(full) );
  QDFZRBS full_pulse_reg ( .D(N162), .TD(full_delay), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(full_pulse) );
  QDFZRBS ptr_reg_1 ( .D(n56), .TD(ptr[0]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[1]) );
  QDFZRBS wr_ptr_reg ( .D(n55), .TD(N4), .SEL(test_se), .CK(hclk), .RB(hresetn), .Q(test_so) );
  QDFZRBS rd_ptr_reg ( .D(n57), .TD(ptr[1]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(N4) );
  QDFZRBS ptr_reg_0 ( .D(n58), .TD(full), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[0]) );
  QDFZRBS fifo_mem_reg_1_31 ( .D(N135), .TD(q_all[62]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[63]) );
  QDFZRBS fifo_mem_reg_1_30 ( .D(N133), .TD(q_all[61]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[62]) );
  QDFZRBS fifo_mem_reg_1_29 ( .D(N131), .TD(q_all[60]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[61]) );
  QDFZRBS fifo_mem_reg_1_28 ( .D(N129), .TD(q_all[59]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[60]) );
  QDFZRBS fifo_mem_reg_1_27 ( .D(N127), .TD(q_all[58]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[59]) );
  QDFZRBS fifo_mem_reg_1_26 ( .D(N125), .TD(q_all[57]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[58]) );
  QDFZRBS fifo_mem_reg_1_25 ( .D(N123), .TD(q_all[56]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[57]) );
  QDFZRBS fifo_mem_reg_1_24 ( .D(N121), .TD(q_all[55]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[56]) );
  QDFZRBS fifo_mem_reg_1_23 ( .D(N119), .TD(q_all[54]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[55]) );
  QDFZRBS fifo_mem_reg_1_22 ( .D(N117), .TD(q_all[53]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[54]) );
  QDFZRBS fifo_mem_reg_1_21 ( .D(N115), .TD(q_all[52]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[53]) );
  QDFZRBS fifo_mem_reg_1_20 ( .D(N113), .TD(q_all[51]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[52]) );
  QDFZRBS fifo_mem_reg_1_19 ( .D(N111), .TD(q_all[50]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[51]) );
  QDFZRBS fifo_mem_reg_1_18 ( .D(N109), .TD(q_all[49]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[50]) );
  QDFZRBS fifo_mem_reg_1_17 ( .D(N107), .TD(q_all[48]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[49]) );
  QDFZRBS fifo_mem_reg_1_16 ( .D(N105), .TD(q_all[47]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[48]) );
  QDFZRBS fifo_mem_reg_1_15 ( .D(N103), .TD(q_all[46]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[47]) );
  QDFZRBS fifo_mem_reg_1_14 ( .D(N101), .TD(q_all[45]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[46]) );
  QDFZRBS fifo_mem_reg_1_13 ( .D(N99), .TD(q_all[44]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[45]) );
  QDFZRBS fifo_mem_reg_1_12 ( .D(N97), .TD(q_all[43]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[44]) );
  QDFZRBS fifo_mem_reg_1_11 ( .D(N95), .TD(q_all[42]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[43]) );
  QDFZRBS fifo_mem_reg_1_10 ( .D(N93), .TD(q_all[41]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[42]) );
  QDFZRBS fifo_mem_reg_1_9 ( .D(N91), .TD(q_all[40]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[41]) );
  QDFZRBS fifo_mem_reg_1_8 ( .D(N89), .TD(q_all[39]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[40]) );
  QDFZRBS fifo_mem_reg_1_7 ( .D(N87), .TD(q_all[38]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[39]) );
  QDFZRBS fifo_mem_reg_1_6 ( .D(N85), .TD(q_all[37]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[38]) );
  QDFZRBS fifo_mem_reg_1_5 ( .D(N83), .TD(q_all[36]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[37]) );
  QDFZRBS fifo_mem_reg_1_4 ( .D(N81), .TD(q_all[35]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[36]) );
  QDFZRBS fifo_mem_reg_1_3 ( .D(N79), .TD(q_all[34]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[35]) );
  QDFZRBS fifo_mem_reg_1_2 ( .D(N77), .TD(q_all[33]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[34]) );
  QDFZRBS fifo_mem_reg_1_1 ( .D(N75), .TD(q_all[32]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[33]) );
  QDFZRBS fifo_mem_reg_1_0 ( .D(N73), .TD(q_all[31]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N134_0_0), .RB(POR), .Q(q_all[32]) );
  QDFZRBS fifo_mem_reg_0_31 ( .D(N71), .TD(q_all[30]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[31]) );
  QDFZRBS fifo_mem_reg_0_30 ( .D(N69), .TD(q_all[29]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[30]) );
  QDFZRBS fifo_mem_reg_0_29 ( .D(N67), .TD(q_all[28]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[29]) );
  QDFZRBS fifo_mem_reg_0_28 ( .D(N65), .TD(q_all[27]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[28]) );
  QDFZRBS fifo_mem_reg_0_27 ( .D(N63), .TD(q_all[26]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[27]) );
  QDFZRBS fifo_mem_reg_0_26 ( .D(N61), .TD(q_all[25]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[26]) );
  QDFZRBS fifo_mem_reg_0_25 ( .D(N59), .TD(q_all[24]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[25]) );
  QDFZRBS fifo_mem_reg_0_24 ( .D(N57), .TD(q_all[23]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[24]) );
  QDFZRBS fifo_mem_reg_0_23 ( .D(N55), .TD(q_all[22]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[23]) );
  QDFZRBS fifo_mem_reg_0_22 ( .D(N53), .TD(q_all[21]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[22]) );
  QDFZRBS fifo_mem_reg_0_21 ( .D(N51), .TD(q_all[20]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[21]) );
  QDFZRBS fifo_mem_reg_0_20 ( .D(N49), .TD(q_all[19]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[20]) );
  QDFZRBS fifo_mem_reg_0_19 ( .D(N47), .TD(q_all[18]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[19]) );
  QDFZRBS fifo_mem_reg_0_18 ( .D(N45), .TD(q_all[17]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[18]) );
  QDFZRBS fifo_mem_reg_0_17 ( .D(N43), .TD(q_all[16]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[17]) );
  QDFZRBS fifo_mem_reg_0_16 ( .D(N41), .TD(q_all[15]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[16]) );
  QDFZRBS fifo_mem_reg_0_15 ( .D(N39), .TD(q_all[14]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[15]) );
  QDFZRBS fifo_mem_reg_0_14 ( .D(N37), .TD(q_all[13]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[14]) );
  QDFZRBS fifo_mem_reg_0_13 ( .D(N35), .TD(q_all[12]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[13]) );
  QDFZRBS fifo_mem_reg_0_12 ( .D(N33), .TD(q_all[11]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[12]) );
  QDFZRBS fifo_mem_reg_0_11 ( .D(N31), .TD(q_all[10]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[11]) );
  QDFZRBS fifo_mem_reg_0_10 ( .D(N29), .TD(q_all[9]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[10]) );
  QDFZRBS fifo_mem_reg_0_9 ( .D(N27), .TD(q_all[8]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[9]) );
  QDFZRBS fifo_mem_reg_0_8 ( .D(N25), .TD(q_all[7]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[8]) );
  QDFZRBS fifo_mem_reg_0_7 ( .D(N23), .TD(q_all[6]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[7]) );
  QDFZRBS fifo_mem_reg_0_6 ( .D(N21), .TD(q_all[5]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[6]) );
  QDFZRBS fifo_mem_reg_0_5 ( .D(N19), .TD(q_all[4]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[5]) );
  QDFZRBS fifo_mem_reg_0_4 ( .D(N17), .TD(q_all[3]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[4]) );
  QDFZRBS fifo_mem_reg_0_3 ( .D(N15), .TD(q_all[2]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[3]) );
  QDFZRBS fifo_mem_reg_0_2 ( .D(N13), .TD(q_all[1]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[2]) );
  QDFZRBS fifo_mem_reg_0_1 ( .D(N11), .TD(q_all[0]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[1]) );
  QDFZRBS fifo_mem_reg_0_0 ( .D(N9), .TD(n78), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N70_0_0), .RB(POR), .Q(q_all[0]) );
endmodule


module des_iv ( hclk, POR, hresetn, clrptr, wr, deswr, data, data_all, q_all, 
        test_mode, test_se, test_si1, test_si2, test_so2, test_so1 );
  input [31:0] data;
  input [63:0] data_all;
  output [63:0] q_all;
  input hclk, POR, hresetn, clrptr, wr, deswr, test_mode, test_se, test_si1,
         test_si2;
  output test_so2, test_so1;
  wire   N5, N7, N9, N11, N13, N15, N17, N19, N21, N23, N25, N27, N29, N31,
         N33, N35, N37, N39, N41, N43, N45, N47, N49, N51, N53, N55, N57, N59,
         N61, N63, N65, N66, N67, N69, N71, N73, N75, N77, N79, N81, N83, N85,
         N87, N89, N91, N93, N95, N97, N99, N101, N103, N105, N107, N109, N111,
         N113, N115, N117, N119, N121, N123, N125, N127, N129, N130, N131,
         CLKGATING_hclk_POWERGATING_hclk_N130_0_0, net1850,
         CLKGATING_hclk_POWERGATING_hclk_N66_0_0, net1855, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n1, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n63;
  wire   [1:0] ptr;

  POWERMODULE_HIGH_des_iv_0_1 POWERGATING_hclk_N130_0 ( .CLK(hclk), .EN(N130), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .TE(n59), .ENOBS(
        net1850) );
  POWERMODULE_HIGH_des_iv_0_0 POWERGATING_hclk_N66_0 ( .CLK(hclk), .EN(N66), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .TE(n59), .ENOBS(
        net1855) );
  SNPS_CLOCK_GATE_OBS_des_iv clk_gate_obs ( .TE(n59), .net1850(net1850), 
        .net1855(net1855), .hclk(hclk), .test_se(test_se), .test_si(test_si2), 
        .test_so(n63) );
  BUF1 U3 ( .I(test_mode), .O(n59) );
  BUF2 U4 ( .I(n7), .O(n51) );
  BUF1 U5 ( .I(n9), .O(n50) );
  BUF2 U6 ( .I(n9), .O(n49) );
  BUF2 U7 ( .I(n9), .O(n1) );
  BUF2 U8 ( .I(n9), .O(n45) );
  BUF2 U9 ( .I(n9), .O(n46) );
  BUF2 U10 ( .I(n9), .O(n47) );
  BUF2 U11 ( .I(n9), .O(n48) );
  BUF1 U12 ( .I(n7), .O(n58) );
  BUF2 U13 ( .I(n7), .O(n57) );
  BUF2 U14 ( .I(n7), .O(n52) );
  BUF2 U15 ( .I(n7), .O(n53) );
  BUF2 U16 ( .I(n7), .O(n54) );
  BUF2 U17 ( .I(n7), .O(n55) );
  BUF2 U18 ( .I(n7), .O(n56) );
  INV2 U19 ( .I(wr), .O(n7) );
  INV2 U20 ( .I(n26), .O(n9) );
  INV2 U21 ( .I(clrptr), .O(n3) );
  ND2 U22 ( .I1(deswr), .I2(n51), .O(n26) );
  AO12 U23 ( .B1(wr), .B2(test_so1), .A1(n50), .O(N130) );
  OAI12S U24 ( .B1(test_so1), .B2(n51), .A1(n26), .O(N66) );
  NR2 U25 ( .I1(n2), .I2(n3), .O(n42) );
  XOR2 U26 ( .I1(n4), .I2(test_so1), .O(n2) );
  NR2 U27 ( .I1(n6), .I2(n3), .O(n44) );
  XOR2 U28 ( .I1(n4), .I2(ptr[0]), .O(n6) );
  MOAI1 U29 ( .A1(n51), .A2(n41), .B1(data_all[48]), .B2(n47), .O(N101) );
  MOAI1 U30 ( .A1(n51), .A2(n40), .B1(data_all[49]), .B2(n1), .O(N103) );
  MOAI1 U31 ( .A1(n51), .A2(n38), .B1(data_all[51]), .B2(n1), .O(N107) );
  MOAI1 U32 ( .A1(n51), .A2(n37), .B1(data_all[52]), .B2(n1), .O(N109) );
  MOAI1 U33 ( .A1(n51), .A2(n36), .B1(data_all[53]), .B2(n1), .O(N111) );
  MOAI1 U34 ( .A1(n51), .A2(n35), .B1(data_all[54]), .B2(n1), .O(N113) );
  MOAI1 U35 ( .A1(n51), .A2(n22), .B1(data_all[3]), .B2(n1), .O(N11) );
  MOAI1 U36 ( .A1(n56), .A2(n24), .B1(data_all[32]), .B2(n48), .O(N69) );
  MOAI1 U37 ( .A1(n56), .A2(n23), .B1(data_all[33]), .B2(n48), .O(N71) );
  MOAI1 U38 ( .A1(n56), .A2(n14), .B1(data_all[34]), .B2(n49), .O(N73) );
  MOAI1 U39 ( .A1(n56), .A2(n22), .B1(data_all[35]), .B2(n49), .O(N75) );
  MOAI1 U40 ( .A1(n56), .A2(n21), .B1(data_all[36]), .B2(n49), .O(N77) );
  MOAI1 U41 ( .A1(n57), .A2(n20), .B1(data_all[37]), .B2(n49), .O(N79) );
  MOAI1 U42 ( .A1(n57), .A2(n19), .B1(data_all[38]), .B2(n49), .O(N81) );
  MOAI1 U43 ( .A1(n57), .A2(n18), .B1(data_all[39]), .B2(n49), .O(N83) );
  MOAI1 U44 ( .A1(n57), .A2(n17), .B1(data_all[40]), .B2(n49), .O(N85) );
  MOAI1 U45 ( .A1(n57), .A2(n16), .B1(data_all[41]), .B2(n49), .O(N87) );
  MOAI1 U46 ( .A1(n57), .A2(n15), .B1(data_all[42]), .B2(n49), .O(N89) );
  MOAI1 U47 ( .A1(n57), .A2(n13), .B1(data_all[43]), .B2(n50), .O(N91) );
  MOAI1 U48 ( .A1(n57), .A2(n12), .B1(data_all[44]), .B2(n50), .O(N93) );
  MOAI1 U49 ( .A1(n52), .A2(n39), .B1(data_all[50]), .B2(n1), .O(N105) );
  MOAI1 U50 ( .A1(n52), .A2(n34), .B1(data_all[55]), .B2(n1), .O(N115) );
  MOAI1 U51 ( .A1(n52), .A2(n33), .B1(data_all[56]), .B2(n1), .O(N117) );
  MOAI1 U52 ( .A1(n52), .A2(n32), .B1(data_all[57]), .B2(n45), .O(N119) );
  MOAI1 U53 ( .A1(n52), .A2(n31), .B1(data_all[58]), .B2(n45), .O(N121) );
  MOAI1 U54 ( .A1(n52), .A2(n30), .B1(data_all[59]), .B2(n45), .O(N123) );
  MOAI1 U55 ( .A1(n52), .A2(n29), .B1(data_all[60]), .B2(n45), .O(N125) );
  MOAI1 U56 ( .A1(n53), .A2(n28), .B1(data_all[61]), .B2(n45), .O(N127) );
  MOAI1 U57 ( .A1(n54), .A2(n27), .B1(data_all[62]), .B2(n45), .O(N129) );
  MOAI1 U58 ( .A1(n52), .A2(n25), .B1(data_all[63]), .B2(n45), .O(N131) );
  MOAI1 U59 ( .A1(n55), .A2(n24), .B1(data_all[0]), .B2(n47), .O(N5) );
  MOAI1 U60 ( .A1(n56), .A2(n23), .B1(data_all[1]), .B2(n48), .O(N7) );
  MOAI1 U61 ( .A1(n57), .A2(n14), .B1(data_all[2]), .B2(n49), .O(N9) );
  MOAI1 U62 ( .A1(n52), .A2(n21), .B1(data_all[4]), .B2(n45), .O(N13) );
  MOAI1 U63 ( .A1(n53), .A2(n20), .B1(data_all[5]), .B2(n45), .O(N15) );
  MOAI1 U64 ( .A1(n53), .A2(n19), .B1(data_all[6]), .B2(n45), .O(N17) );
  MOAI1 U65 ( .A1(n53), .A2(n18), .B1(data_all[7]), .B2(n46), .O(N19) );
  MOAI1 U66 ( .A1(n53), .A2(n17), .B1(data_all[8]), .B2(n46), .O(N21) );
  MOAI1 U67 ( .A1(n53), .A2(n16), .B1(data_all[9]), .B2(n46), .O(N23) );
  MOAI1 U68 ( .A1(n53), .A2(n15), .B1(data_all[10]), .B2(n46), .O(N25) );
  MOAI1 U69 ( .A1(n53), .A2(n13), .B1(data_all[11]), .B2(n46), .O(N27) );
  MOAI1 U70 ( .A1(n53), .A2(n12), .B1(data_all[12]), .B2(n46), .O(N29) );
  MOAI1 U71 ( .A1(n54), .A2(n11), .B1(data_all[13]), .B2(n46), .O(N31) );
  MOAI1 U72 ( .A1(n54), .A2(n10), .B1(data_all[14]), .B2(n46), .O(N33) );
  MOAI1 U73 ( .A1(n54), .A2(n8), .B1(data_all[15]), .B2(n46), .O(N35) );
  MOAI1 U74 ( .A1(n54), .A2(n41), .B1(data_all[16]), .B2(n46), .O(N37) );
  MOAI1 U75 ( .A1(n54), .A2(n40), .B1(data_all[17]), .B2(n47), .O(N39) );
  MOAI1 U76 ( .A1(n54), .A2(n39), .B1(data_all[18]), .B2(n47), .O(N41) );
  MOAI1 U77 ( .A1(n54), .A2(n38), .B1(data_all[19]), .B2(n47), .O(N43) );
  MOAI1 U78 ( .A1(n54), .A2(n37), .B1(data_all[20]), .B2(n47), .O(N45) );
  MOAI1 U79 ( .A1(n55), .A2(n36), .B1(data_all[21]), .B2(n47), .O(N47) );
  MOAI1 U80 ( .A1(n55), .A2(n35), .B1(data_all[22]), .B2(n47), .O(N49) );
  MOAI1 U81 ( .A1(n55), .A2(n34), .B1(data_all[23]), .B2(n47), .O(N51) );
  MOAI1 U82 ( .A1(n55), .A2(n33), .B1(data_all[24]), .B2(n47), .O(N53) );
  MOAI1 U83 ( .A1(n55), .A2(n32), .B1(data_all[25]), .B2(n48), .O(N55) );
  MOAI1 U84 ( .A1(n55), .A2(n31), .B1(data_all[26]), .B2(n48), .O(N57) );
  MOAI1 U85 ( .A1(n55), .A2(n30), .B1(data_all[27]), .B2(n48), .O(N59) );
  MOAI1 U86 ( .A1(n55), .A2(n29), .B1(data_all[28]), .B2(n48), .O(N61) );
  MOAI1 U87 ( .A1(n56), .A2(n28), .B1(data_all[29]), .B2(n48), .O(N63) );
  MOAI1 U88 ( .A1(n56), .A2(n27), .B1(data_all[30]), .B2(n48), .O(N65) );
  MOAI1 U89 ( .A1(n56), .A2(n25), .B1(data_all[31]), .B2(n48), .O(N67) );
  MOAI1 U90 ( .A1(n58), .A2(n11), .B1(data_all[45]), .B2(n50), .O(N95) );
  MOAI1 U91 ( .A1(n58), .A2(n10), .B1(data_all[46]), .B2(n50), .O(N97) );
  MOAI1 U92 ( .A1(n58), .A2(n8), .B1(data_all[47]), .B2(n1), .O(N99) );
  OR2 U93 ( .I1(n58), .I2(ptr[1]), .O(n4) );
  INV2 U94 ( .I(data[1]), .O(n23) );
  INV2 U95 ( .I(data[2]), .O(n14) );
  INV2 U96 ( .I(data[3]), .O(n22) );
  INV2 U97 ( .I(data[4]), .O(n21) );
  INV2 U98 ( .I(data[5]), .O(n20) );
  INV2 U99 ( .I(data[6]), .O(n19) );
  INV2 U100 ( .I(data[7]), .O(n18) );
  INV2 U101 ( .I(data[9]), .O(n16) );
  INV2 U102 ( .I(data[10]), .O(n15) );
  INV2 U103 ( .I(data[11]), .O(n13) );
  INV2 U104 ( .I(data[12]), .O(n12) );
  INV2 U105 ( .I(data[13]), .O(n11) );
  INV2 U106 ( .I(data[14]), .O(n10) );
  INV2 U107 ( .I(data[15]), .O(n8) );
  INV2 U108 ( .I(data[17]), .O(n40) );
  INV2 U109 ( .I(data[18]), .O(n39) );
  INV2 U110 ( .I(data[19]), .O(n38) );
  INV2 U111 ( .I(data[20]), .O(n37) );
  INV2 U112 ( .I(data[21]), .O(n36) );
  INV2 U113 ( .I(data[22]), .O(n35) );
  INV2 U114 ( .I(data[23]), .O(n34) );
  INV2 U115 ( .I(data[25]), .O(n32) );
  INV2 U116 ( .I(data[26]), .O(n31) );
  INV2 U117 ( .I(data[27]), .O(n30) );
  INV2 U118 ( .I(data[28]), .O(n29) );
  INV2 U119 ( .I(data[29]), .O(n28) );
  INV2 U120 ( .I(data[30]), .O(n27) );
  INV2 U121 ( .I(data[31]), .O(n25) );
  INV2 U122 ( .I(data[0]), .O(n24) );
  INV2 U123 ( .I(data[8]), .O(n17) );
  INV2 U124 ( .I(data[16]), .O(n41) );
  INV2 U125 ( .I(data[24]), .O(n33) );
  NR2 U126 ( .I1(n5), .I2(n3), .O(n43) );
  AOI12S U127 ( .B1(ptr[0]), .B2(wr), .A1(ptr[1]), .O(n5) );
  QDFZRBS ptr_reg_1 ( .D(n43), .TD(ptr[0]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[1]) );
  QDFZRBS ptr_reg_0 ( .D(n44), .TD(q_all[63]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[0]) );
  QDFZRBS fifo_mem_reg_0_30 ( .D(N65), .TD(q_all[29]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[30]) );
  QDFZRBS fifo_mem_reg_0_28 ( .D(N61), .TD(q_all[27]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[28]) );
  QDFZRBS fifo_mem_reg_0_26 ( .D(N57), .TD(q_all[25]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[26]) );
  QDFZRBS fifo_mem_reg_0_24 ( .D(N53), .TD(q_all[23]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[24]) );
  QDFZRBS fifo_mem_reg_0_22 ( .D(N49), .TD(q_all[21]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[22]) );
  QDFZRBS fifo_mem_reg_0_20 ( .D(N45), .TD(q_all[19]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[20]) );
  QDFZRBS fifo_mem_reg_0_18 ( .D(N41), .TD(q_all[17]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[18]) );
  QDFZRBS fifo_mem_reg_0_16 ( .D(N37), .TD(q_all[15]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[16]) );
  QDFZRBS fifo_mem_reg_0_14 ( .D(N33), .TD(q_all[13]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[14]) );
  QDFZRBS fifo_mem_reg_0_12 ( .D(N29), .TD(q_all[11]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[12]) );
  QDFZRBS fifo_mem_reg_0_10 ( .D(N25), .TD(q_all[9]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[10]) );
  QDFZRBS fifo_mem_reg_0_8 ( .D(N21), .TD(q_all[7]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[8]) );
  QDFZRBS fifo_mem_reg_0_6 ( .D(N17), .TD(q_all[5]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[6]) );
  QDFZRBS fifo_mem_reg_0_4 ( .D(N13), .TD(q_all[3]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[4]) );
  QDFZRBS fifo_mem_reg_0_2 ( .D(N9), .TD(q_all[1]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[2]) );
  QDFZRBS fifo_mem_reg_0_0 ( .D(N5), .TD(n63), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[0]) );
  QDFZRBS fifo_mem_reg_1_30 ( .D(N129), .TD(q_all[61]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[62]) );
  QDFZRBS fifo_mem_reg_1_28 ( .D(N125), .TD(q_all[59]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[60]) );
  QDFZRBS fifo_mem_reg_1_26 ( .D(N121), .TD(q_all[57]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[58]) );
  QDFZRBS fifo_mem_reg_1_24 ( .D(N117), .TD(q_all[55]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[56]) );
  QDFZRBS fifo_mem_reg_1_22 ( .D(N113), .TD(q_all[53]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[54]) );
  QDFZRBS fifo_mem_reg_1_20 ( .D(N109), .TD(q_all[51]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[52]) );
  QDFZRBS fifo_mem_reg_1_18 ( .D(N105), .TD(q_all[49]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[50]) );
  QDFZRBS fifo_mem_reg_1_16 ( .D(N101), .TD(q_all[47]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[48]) );
  QDFZRBS fifo_mem_reg_1_14 ( .D(N97), .TD(q_all[45]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[46]) );
  QDFZRBS fifo_mem_reg_1_12 ( .D(N93), .TD(q_all[43]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[44]) );
  QDFZRBS fifo_mem_reg_1_10 ( .D(N89), .TD(q_all[41]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[42]) );
  QDFZRBS fifo_mem_reg_1_8 ( .D(N85), .TD(q_all[39]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[40]) );
  QDFZRBS fifo_mem_reg_1_6 ( .D(N81), .TD(q_all[37]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[38]) );
  QDFZRBS fifo_mem_reg_1_4 ( .D(N77), .TD(q_all[35]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[36]) );
  QDFZRBS fifo_mem_reg_1_2 ( .D(N73), .TD(q_all[33]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[34]) );
  QDFZRBS fifo_mem_reg_1_0 ( .D(N69), .TD(q_all[31]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[32]) );
  QDFZRBS fifo_mem_reg_0_15 ( .D(N35), .TD(q_all[14]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[15]) );
  QDFZRBS fifo_mem_reg_1_23 ( .D(N115), .TD(q_all[54]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[55]) );
  QDFZRBS fifo_mem_reg_1_13 ( .D(N95), .TD(q_all[44]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[45]) );
  QDFZRBS fifo_mem_reg_1_11 ( .D(N91), .TD(q_all[42]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[43]) );
  QDFZRBS fifo_mem_reg_1_9 ( .D(N87), .TD(q_all[40]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[41]) );
  QDFZRBS fifo_mem_reg_0_31 ( .D(N67), .TD(q_all[30]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[31]) );
  QDFZRBS fifo_mem_reg_0_29 ( .D(N63), .TD(test_si1), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[29]) );
  QDFZRBS fifo_mem_reg_0_27 ( .D(N59), .TD(q_all[26]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[27]) );
  QDFZRBS fifo_mem_reg_0_25 ( .D(N55), .TD(q_all[24]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[25]) );
  QDFZRBS fifo_mem_reg_0_23 ( .D(N51), .TD(q_all[22]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[23]) );
  QDFZRBS fifo_mem_reg_0_21 ( .D(N47), .TD(q_all[20]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[21]) );
  QDFZRBS fifo_mem_reg_0_19 ( .D(N43), .TD(q_all[18]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[19]) );
  QDFZRBS fifo_mem_reg_0_17 ( .D(N39), .TD(q_all[16]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[17]) );
  QDFZRBS fifo_mem_reg_0_13 ( .D(N31), .TD(q_all[12]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[13]) );
  QDFZRBS fifo_mem_reg_0_11 ( .D(N27), .TD(q_all[10]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[11]) );
  QDFZRBS fifo_mem_reg_0_9 ( .D(N23), .TD(q_all[8]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[9]) );
  QDFZRBS fifo_mem_reg_0_7 ( .D(N19), .TD(q_all[6]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[7]) );
  QDFZRBS fifo_mem_reg_0_5 ( .D(N15), .TD(q_all[4]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[5]) );
  QDFZRBS fifo_mem_reg_0_3 ( .D(N11), .TD(q_all[2]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[3]) );
  QDFZRBS fifo_mem_reg_0_1 ( .D(N7), .TD(q_all[0]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .RB(POR), .Q(q_all[1]) );
  QDFZRBS fifo_mem_reg_1_29 ( .D(N127), .TD(q_all[60]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[61]) );
  QDFZRBS fifo_mem_reg_1_27 ( .D(N123), .TD(q_all[58]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[59]) );
  QDFZRBS fifo_mem_reg_1_25 ( .D(N119), .TD(q_all[56]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[57]) );
  QDFZRBS fifo_mem_reg_1_21 ( .D(N111), .TD(q_all[52]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[53]) );
  QDFZRBS fifo_mem_reg_1_19 ( .D(N107), .TD(q_all[50]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[51]) );
  QDFZRBS fifo_mem_reg_1_17 ( .D(N103), .TD(q_all[48]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[49]) );
  QDFZRBS fifo_mem_reg_1_15 ( .D(N99), .TD(q_all[46]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[47]) );
  QDFZRBS fifo_mem_reg_1_7 ( .D(N83), .TD(q_all[38]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[39]) );
  QDFZRBS fifo_mem_reg_1_5 ( .D(N79), .TD(q_all[36]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[37]) );
  QDFZRBS fifo_mem_reg_1_3 ( .D(N75), .TD(q_all[34]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[35]) );
  QDFZRBS fifo_mem_reg_1_1 ( .D(N71), .TD(q_all[32]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[33]) );
  QDFZRBS fifo_mem_reg_1_31 ( .D(N131), .TD(q_all[62]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N130_0_0), .RB(POR), .Q(q_all[63]) );
  QDFZRBS wr_ptr_reg ( .D(n42), .TD(ptr[1]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(test_so1) );
  QDBHN LOCKUP ( .CKB(CLKGATING_hclk_POWERGATING_hclk_N66_0_0), .D(q_all[28]), 
        .Q(test_so2) );
endmodule


module des_key ( hresetn, clrptr, hclk, wr, data, q1_all, q2_all, q3_all, 
        test_mode, test_se, test_si1, test_si2, test_so2, test_so1 );
  input [31:0] data;
  output [63:0] q1_all;
  output [63:0] q2_all;
  output [63:0] q3_all;
  input hresetn, clrptr, hclk, wr, test_mode, test_se, test_si1, test_si2;
  output test_so2, test_so1;
  wire   N83, N115, N147, N179, N211, N243,
         CLKGATING_hclk_POWERGATING_hclk_N243_0_0, net1889,
         CLKGATING_hclk_POWERGATING_hclk_N211_0_0, net1894,
         CLKGATING_hclk_POWERGATING_hclk_N179_0_0, net1899,
         CLKGATING_hclk_POWERGATING_hclk_N147_0_0, net1904,
         CLKGATING_hclk_POWERGATING_hclk_N115_0_0, net1909,
         CLKGATING_hclk_POWERGATING_hclk_N83_0_0, net1914, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n2, n59, n60, wr_ptr_1_, wr_ptr_0_, n5;
  wire   [2:0] ptr;

  POWERMODULE_HIGH_des_key_0_5 POWERGATING_hclk_N243_0 ( .CLK(hclk), .EN(N243), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .TE(n60), .ENOBS(
        net1889) );
  POWERMODULE_HIGH_des_key_0_4 POWERGATING_hclk_N211_0 ( .CLK(hclk), .EN(N211), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .TE(n59), .ENOBS(
        net1894) );
  POWERMODULE_HIGH_des_key_0_3 POWERGATING_hclk_N179_0 ( .CLK(hclk), .EN(N179), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .TE(n60), .ENOBS(
        net1899) );
  POWERMODULE_HIGH_des_key_0_2 POWERGATING_hclk_N147_0 ( .CLK(hclk), .EN(N147), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .TE(n60), .ENOBS(
        net1904) );
  POWERMODULE_HIGH_des_key_0_1 POWERGATING_hclk_N115_0 ( .CLK(hclk), .EN(N115), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .TE(n59), .ENOBS(
        net1909) );
  POWERMODULE_HIGH_des_key_0_0 POWERGATING_hclk_N83_0 ( .CLK(hclk), .EN(N83), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .TE(n59), .ENOBS(
        net1914) );
  SNPS_CLOCK_GATE_OBS_des_key clk_gate_obs ( .TE(n59), .net1889(net1889), 
        .net1894(net1894), .net1899(net1899), .net1904(net1904), .net1909(
        net1909), .net1914(net1914), .hclk(hclk), .test_se(test_se), .test_si(
        test_si2), .test_so(n5) );
  TIE1 U3 ( .O(n2) );
  INV2 U4 ( .I(n2), .O(q3_all[0]) );
  INV2 U5 ( .I(n2), .O(q3_all[8]) );
  INV2 U6 ( .I(n2), .O(q3_all[16]) );
  INV2 U7 ( .I(n2), .O(q3_all[24]) );
  INV2 U8 ( .I(n2), .O(q3_all[32]) );
  INV2 U9 ( .I(n2), .O(q3_all[40]) );
  INV2 U10 ( .I(n2), .O(q3_all[48]) );
  INV2 U11 ( .I(n2), .O(q3_all[56]) );
  INV2 U12 ( .I(n2), .O(q2_all[0]) );
  INV2 U13 ( .I(n2), .O(q2_all[8]) );
  INV2 U14 ( .I(n2), .O(q2_all[16]) );
  INV2 U15 ( .I(n2), .O(q2_all[24]) );
  INV2 U16 ( .I(n2), .O(q2_all[32]) );
  INV2 U17 ( .I(n2), .O(q2_all[40]) );
  INV2 U18 ( .I(n2), .O(q2_all[48]) );
  INV2 U19 ( .I(n2), .O(q2_all[56]) );
  INV2 U20 ( .I(n2), .O(q1_all[0]) );
  INV2 U21 ( .I(n2), .O(q1_all[8]) );
  INV2 U22 ( .I(n2), .O(q1_all[16]) );
  INV2 U23 ( .I(n2), .O(q1_all[24]) );
  INV2 U24 ( .I(n2), .O(q1_all[32]) );
  INV2 U25 ( .I(n2), .O(q1_all[40]) );
  INV2 U26 ( .I(n2), .O(q1_all[48]) );
  INV2 U27 ( .I(n2), .O(q1_all[56]) );
  ND2 U28 ( .I1(n27), .I2(n11), .O(n28) );
  INV2 U29 ( .I(wr_ptr_1_), .O(n19) );
  ND3 U30 ( .I1(wr_ptr_1_), .I2(clrptr), .I3(test_so1), .O(n13) );
  NR2 U31 ( .I1(n28), .I2(n36), .O(N83) );
  NR2P U32 ( .I1(n28), .I2(n26), .O(n22) );
  NR3P U33 ( .I1(n21), .I2(n19), .I3(n35), .O(N179) );
  NR3P U34 ( .I1(n28), .I2(n19), .I3(n35), .O(N147) );
  NR3P U35 ( .I1(n36), .I2(n11), .I3(n27), .O(N243) );
  ND2P U36 ( .I1(wr), .I2(n19), .O(n36) );
  INV2 U37 ( .I(wr), .O(n35) );
  NR2 U38 ( .I1(n21), .I2(n36), .O(N115) );
  INV2 U39 ( .I(n14), .O(n26) );
  ND2P U40 ( .I1(clrptr), .I2(n26), .O(n17) );
  ND3 U41 ( .I1(n27), .I2(n19), .I3(n14), .O(n16) );
  OAI112S U42 ( .C1(n18), .C2(n19), .A1(n20), .B1(n13), .O(n38) );
  ND3 U43 ( .I1(n14), .I2(n19), .I3(n15), .O(n20) );
  NR2 U44 ( .I1(n22), .I2(n23), .O(n18) );
  INV2 U45 ( .I(n17), .O(n23) );
  MOAI1 U46 ( .A1(n32), .A2(n17), .B1(n14), .B2(n32), .O(n42) );
  INV2 U47 ( .I(clrptr), .O(n29) );
  INV2 U48 ( .I(n21), .O(n15) );
  NR3P U49 ( .I1(n36), .I2(wr_ptr_0_), .I3(n11), .O(N211) );
  ND2P U50 ( .I1(wr_ptr_0_), .I2(n11), .O(n21) );
  INV2 U51 ( .I(wr_ptr_0_), .O(n27) );
  AOI112P U52 ( .C1(ptr[1]), .C2(ptr[2]), .A1(n29), .B1(n35), .O(n14) );
  OAI12S U53 ( .B1(n29), .B2(n30), .A1(n31), .O(n40) );
  INV2 U54 ( .I(ptr[2]), .O(n30) );
  ND3 U55 ( .I1(n14), .I2(ptr[1]), .I3(ptr[0]), .O(n31) );
  OAI112S U56 ( .C1(n10), .C2(n11), .A1(n12), .B1(n13), .O(n37) );
  ND3 U57 ( .I1(n14), .I2(wr_ptr_1_), .I3(n15), .O(n12) );
  AN2 U58 ( .I1(n16), .I2(n17), .O(n10) );
  MOAI1 U59 ( .A1(n32), .A2(n33), .B1(ptr[1]), .B2(n34), .O(n41) );
  OR2 U60 ( .I1(n26), .I2(ptr[1]), .O(n33) );
  OAI12S U61 ( .B1(ptr[0]), .B2(n26), .A1(n17), .O(n34) );
  OR3B2 U62 ( .I1(n22), .B1(n16), .B2(n24), .O(n39) );
  OAI112S U63 ( .C1(n25), .C2(n26), .A1(clrptr), .B1(wr_ptr_0_), .O(n24) );
  NR2 U64 ( .I1(n19), .I2(n11), .O(n25) );
  INV2 U65 ( .I(ptr[0]), .O(n32) );
  BUF1 U66 ( .I(test_mode), .O(n59) );
  BUF1 U67 ( .I(test_mode), .O(n60) );
  QDFZRBS ptr_reg_0 ( .D(n42), .TD(q3_all[63]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[0]) );
  QDFZRBS ptr_reg_2 ( .D(n40), .TD(ptr[1]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[2]) );
  QDFZRBS fifo_mem_reg_3_31 ( .D(data[31]), .TD(q2_all[62]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[63]) );
  QDFZRBS fifo_mem_reg_3_30 ( .D(data[30]), .TD(q2_all[61]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[62]) );
  QDFZRBS fifo_mem_reg_3_29 ( .D(data[29]), .TD(q2_all[60]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[61]) );
  QDFZRBS fifo_mem_reg_3_28 ( .D(data[28]), .TD(q2_all[59]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[60]) );
  QDFZRBS fifo_mem_reg_3_27 ( .D(data[27]), .TD(q2_all[58]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[59]) );
  QDFZRBS fifo_mem_reg_3_26 ( .D(data[26]), .TD(q2_all[57]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[58]) );
  QDFZRBS fifo_mem_reg_3_25 ( .D(data[25]), .TD(q2_all[55]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[57]) );
  QDFZRBS fifo_mem_reg_3_23 ( .D(data[23]), .TD(q2_all[54]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[55]) );
  QDFZRBS fifo_mem_reg_3_22 ( .D(data[22]), .TD(q2_all[53]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[54]) );
  QDFZRBS fifo_mem_reg_3_21 ( .D(data[21]), .TD(q2_all[52]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[53]) );
  QDFZRBS fifo_mem_reg_3_20 ( .D(data[20]), .TD(q2_all[51]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[52]) );
  QDFZRBS fifo_mem_reg_3_19 ( .D(data[19]), .TD(q2_all[50]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[51]) );
  QDFZRBS fifo_mem_reg_3_18 ( .D(data[18]), .TD(q2_all[49]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[50]) );
  QDFZRBS fifo_mem_reg_3_17 ( .D(data[17]), .TD(q2_all[47]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[49]) );
  QDFZRBS fifo_mem_reg_3_15 ( .D(data[15]), .TD(q2_all[46]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[47]) );
  QDFZRBS fifo_mem_reg_3_14 ( .D(data[14]), .TD(q2_all[45]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[46]) );
  QDFZRBS fifo_mem_reg_3_13 ( .D(data[13]), .TD(q2_all[44]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[45]) );
  QDFZRBS fifo_mem_reg_3_12 ( .D(data[12]), .TD(q2_all[43]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[44]) );
  QDFZRBS fifo_mem_reg_3_11 ( .D(data[11]), .TD(q2_all[42]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[43]) );
  QDFZRBS fifo_mem_reg_3_10 ( .D(data[10]), .TD(q2_all[41]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(
        q2_all[42]) );
  QDFZRBS fifo_mem_reg_3_9 ( .D(data[9]), .TD(q2_all[39]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[41]) );
  QDFZRBS fifo_mem_reg_3_7 ( .D(data[7]), .TD(q2_all[38]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[39]) );
  QDFZRBS fifo_mem_reg_3_6 ( .D(data[6]), .TD(q2_all[37]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[38]) );
  QDFZRBS fifo_mem_reg_3_5 ( .D(data[5]), .TD(q2_all[36]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[37]) );
  QDFZRBS fifo_mem_reg_3_4 ( .D(data[4]), .TD(q2_all[35]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[36]) );
  QDFZRBS fifo_mem_reg_3_3 ( .D(data[3]), .TD(q2_all[34]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[35]) );
  QDFZRBS fifo_mem_reg_3_2 ( .D(data[2]), .TD(q2_all[33]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[34]) );
  QDFZRBS fifo_mem_reg_3_1 ( .D(data[1]), .TD(q2_all[31]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N179_0_0), .RB(hresetn), .Q(q2_all[33]) );
  QDFZRBS fifo_mem_reg_2_31 ( .D(data[31]), .TD(q2_all[30]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[31]) );
  QDFZRBS fifo_mem_reg_2_30 ( .D(data[30]), .TD(q2_all[29]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[30]) );
  QDFZRBS fifo_mem_reg_2_29 ( .D(data[29]), .TD(q2_all[28]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[29]) );
  QDFZRBS fifo_mem_reg_2_28 ( .D(data[28]), .TD(q2_all[27]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[28]) );
  QDFZRBS fifo_mem_reg_2_27 ( .D(data[27]), .TD(q2_all[26]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[27]) );
  QDFZRBS fifo_mem_reg_2_26 ( .D(data[26]), .TD(q2_all[25]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[26]) );
  QDFZRBS fifo_mem_reg_2_25 ( .D(data[25]), .TD(q2_all[23]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[25]) );
  QDFZRBS fifo_mem_reg_2_23 ( .D(data[23]), .TD(q2_all[22]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[23]) );
  QDFZRBS fifo_mem_reg_2_22 ( .D(data[22]), .TD(q2_all[21]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[22]) );
  QDFZRBS fifo_mem_reg_2_21 ( .D(data[21]), .TD(q2_all[20]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[21]) );
  QDFZRBS fifo_mem_reg_2_20 ( .D(data[20]), .TD(q2_all[19]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[20]) );
  QDFZRBS fifo_mem_reg_2_19 ( .D(data[19]), .TD(q2_all[18]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[19]) );
  QDFZRBS fifo_mem_reg_2_18 ( .D(data[18]), .TD(q2_all[17]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[18]) );
  QDFZRBS fifo_mem_reg_2_17 ( .D(data[17]), .TD(test_si1), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[17]) );
  QDFZRBS fifo_mem_reg_2_15 ( .D(data[15]), .TD(q2_all[14]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[15]) );
  QDFZRBS fifo_mem_reg_2_14 ( .D(data[14]), .TD(q2_all[13]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[14]) );
  QDFZRBS fifo_mem_reg_2_13 ( .D(data[13]), .TD(q2_all[12]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[13]) );
  QDFZRBS fifo_mem_reg_2_12 ( .D(data[12]), .TD(q2_all[11]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[12]) );
  QDFZRBS fifo_mem_reg_2_11 ( .D(data[11]), .TD(q2_all[10]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[11]) );
  QDFZRBS fifo_mem_reg_2_10 ( .D(data[10]), .TD(q2_all[9]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(
        q2_all[10]) );
  QDFZRBS fifo_mem_reg_2_9 ( .D(data[9]), .TD(q2_all[7]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[9])
         );
  QDFZRBS fifo_mem_reg_2_7 ( .D(data[7]), .TD(q2_all[6]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[7])
         );
  QDFZRBS fifo_mem_reg_2_6 ( .D(data[6]), .TD(q2_all[5]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[6])
         );
  QDFZRBS fifo_mem_reg_2_5 ( .D(data[5]), .TD(q2_all[4]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[5])
         );
  QDFZRBS fifo_mem_reg_2_4 ( .D(data[4]), .TD(q2_all[3]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[4])
         );
  QDFZRBS fifo_mem_reg_2_3 ( .D(data[3]), .TD(q2_all[2]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[3])
         );
  QDFZRBS fifo_mem_reg_2_2 ( .D(data[2]), .TD(q2_all[1]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[2])
         );
  QDFZRBS fifo_mem_reg_2_1 ( .D(data[1]), .TD(q1_all[63]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .RB(hresetn), .Q(q2_all[1])
         );
  QDFZRBS fifo_mem_reg_1_31 ( .D(data[31]), .TD(q1_all[62]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[63]) );
  QDFZRBS fifo_mem_reg_1_28 ( .D(data[28]), .TD(q1_all[59]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[60]) );
  QDFZRBS fifo_mem_reg_1_27 ( .D(data[27]), .TD(q1_all[58]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[59]) );
  QDFZRBS fifo_mem_reg_1_26 ( .D(data[26]), .TD(q1_all[57]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[58]) );
  QDFZRBS fifo_mem_reg_1_25 ( .D(data[25]), .TD(q1_all[55]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[57]) );
  QDFZRBS fifo_mem_reg_1_23 ( .D(data[23]), .TD(q1_all[54]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[55]) );
  QDFZRBS fifo_mem_reg_1_22 ( .D(data[22]), .TD(q1_all[53]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[54]) );
  QDFZRBS fifo_mem_reg_1_21 ( .D(data[21]), .TD(q1_all[52]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[53]) );
  QDFZRBS fifo_mem_reg_1_20 ( .D(data[20]), .TD(q1_all[51]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[52]) );
  QDFZRBS fifo_mem_reg_1_19 ( .D(data[19]), .TD(q1_all[50]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[51]) );
  QDFZRBS fifo_mem_reg_1_18 ( .D(data[18]), .TD(q1_all[49]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[50]) );
  QDFZRBS fifo_mem_reg_1_17 ( .D(data[17]), .TD(q1_all[47]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[49]) );
  QDFZRBS fifo_mem_reg_1_15 ( .D(data[15]), .TD(q1_all[46]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[47]) );
  QDFZRBS fifo_mem_reg_1_13 ( .D(data[13]), .TD(q1_all[44]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[45]) );
  QDFZRBS fifo_mem_reg_1_12 ( .D(data[12]), .TD(q1_all[43]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[44]) );
  QDFZRBS fifo_mem_reg_1_11 ( .D(data[11]), .TD(q1_all[42]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[43]) );
  QDFZRBS fifo_mem_reg_1_10 ( .D(data[10]), .TD(q1_all[41]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[42]) );
  QDFZRBS fifo_mem_reg_1_9 ( .D(data[9]), .TD(q1_all[39]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[41]) );
  QDFZRBS fifo_mem_reg_1_7 ( .D(data[7]), .TD(q1_all[38]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[39]) );
  QDFZRBS fifo_mem_reg_1_6 ( .D(data[6]), .TD(q1_all[37]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[38]) );
  QDFZRBS fifo_mem_reg_1_5 ( .D(data[5]), .TD(q1_all[36]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[37]) );
  QDFZRBS fifo_mem_reg_1_4 ( .D(data[4]), .TD(q1_all[35]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[36]) );
  QDFZRBS fifo_mem_reg_1_3 ( .D(data[3]), .TD(q1_all[34]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[35]) );
  QDFZRBS fifo_mem_reg_1_2 ( .D(data[2]), .TD(q1_all[33]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[34]) );
  QDFZRBS fifo_mem_reg_1_1 ( .D(data[1]), .TD(q1_all[31]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(q1_all[33]) );
  QDFZRBS fifo_mem_reg_0_31 ( .D(data[31]), .TD(q1_all[30]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[31]) );
  QDFZRBS fifo_mem_reg_0_29 ( .D(data[29]), .TD(q1_all[28]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[29]) );
  QDFZRBS fifo_mem_reg_0_28 ( .D(data[28]), .TD(q1_all[27]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[28]) );
  QDFZRBS fifo_mem_reg_0_27 ( .D(data[27]), .TD(q1_all[26]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[27]) );
  QDFZRBS fifo_mem_reg_0_26 ( .D(data[26]), .TD(q1_all[25]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[26]) );
  QDFZRBS fifo_mem_reg_0_25 ( .D(data[25]), .TD(q1_all[23]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[25]) );
  QDFZRBS fifo_mem_reg_0_23 ( .D(data[23]), .TD(q1_all[22]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[23]) );
  QDFZRBS fifo_mem_reg_0_22 ( .D(data[22]), .TD(q1_all[21]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[22]) );
  QDFZRBS fifo_mem_reg_0_20 ( .D(data[20]), .TD(q1_all[19]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[20]) );
  QDFZRBS fifo_mem_reg_0_19 ( .D(data[19]), .TD(q1_all[18]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[19]) );
  QDFZRBS fifo_mem_reg_0_18 ( .D(data[18]), .TD(q1_all[17]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[18]) );
  QDFZRBS fifo_mem_reg_0_17 ( .D(data[17]), .TD(q1_all[15]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[17]) );
  QDFZRBS fifo_mem_reg_0_15 ( .D(data[15]), .TD(q1_all[14]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[15]) );
  QDFZRBS fifo_mem_reg_0_14 ( .D(data[14]), .TD(q1_all[13]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[14]) );
  QDFZRBS fifo_mem_reg_0_11 ( .D(data[11]), .TD(q1_all[10]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[11]) );
  QDFZRBS fifo_mem_reg_0_10 ( .D(data[10]), .TD(q1_all[9]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[10]) );
  QDFZRBS fifo_mem_reg_0_9 ( .D(data[9]), .TD(q1_all[7]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[9])
         );
  QDFZRBS fifo_mem_reg_0_7 ( .D(data[7]), .TD(q1_all[6]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[7])
         );
  QDFZRBS fifo_mem_reg_0_6 ( .D(data[6]), .TD(q1_all[5]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[6])
         );
  QDFZRBS fifo_mem_reg_0_4 ( .D(data[4]), .TD(q1_all[3]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[4])
         );
  QDFZRBS fifo_mem_reg_0_3 ( .D(data[3]), .TD(q1_all[2]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[3])
         );
  QDFZRBS fifo_mem_reg_0_2 ( .D(data[2]), .TD(q1_all[1]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[2])
         );
  QDFZRBS fifo_mem_reg_0_1 ( .D(data[1]), .TD(n5), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[1])
         );
  QDFZRBS fifo_mem_reg_5_31 ( .D(data[31]), .TD(q3_all[62]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[63]) );
  QDFZRBS fifo_mem_reg_5_28 ( .D(data[28]), .TD(q3_all[59]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[60]) );
  QDFZRBS fifo_mem_reg_5_27 ( .D(data[27]), .TD(q3_all[58]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[59]) );
  QDFZRBS fifo_mem_reg_5_26 ( .D(data[26]), .TD(q3_all[57]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[58]) );
  QDFZRBS fifo_mem_reg_5_25 ( .D(data[25]), .TD(q3_all[55]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[57]) );
  QDFZRBS fifo_mem_reg_5_23 ( .D(data[23]), .TD(q3_all[54]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[55]) );
  QDFZRBS fifo_mem_reg_5_21 ( .D(data[21]), .TD(q3_all[52]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[53]) );
  QDFZRBS fifo_mem_reg_5_20 ( .D(data[20]), .TD(q3_all[51]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[52]) );
  QDFZRBS fifo_mem_reg_5_19 ( .D(data[19]), .TD(q3_all[50]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[51]) );
  QDFZRBS fifo_mem_reg_5_18 ( .D(data[18]), .TD(q3_all[49]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[50]) );
  QDFZRBS fifo_mem_reg_5_17 ( .D(data[17]), .TD(q3_all[47]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[49]) );
  QDFZRBS fifo_mem_reg_5_15 ( .D(data[15]), .TD(q3_all[46]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[47]) );
  QDFZRBS fifo_mem_reg_5_12 ( .D(data[12]), .TD(q3_all[43]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[44]) );
  QDFZRBS fifo_mem_reg_5_11 ( .D(data[11]), .TD(q3_all[42]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[43]) );
  QDFZRBS fifo_mem_reg_5_10 ( .D(data[10]), .TD(q3_all[41]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[42]) );
  QDFZRBS fifo_mem_reg_5_9 ( .D(data[9]), .TD(q3_all[39]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[41]) );
  QDFZRBS fifo_mem_reg_5_7 ( .D(data[7]), .TD(q3_all[38]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[39]) );
  QDFZRBS fifo_mem_reg_5_5 ( .D(data[5]), .TD(q3_all[36]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[37]) );
  QDFZRBS fifo_mem_reg_5_4 ( .D(data[4]), .TD(q3_all[35]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[36]) );
  QDFZRBS fifo_mem_reg_5_3 ( .D(data[3]), .TD(q3_all[34]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[35]) );
  QDFZRBS fifo_mem_reg_5_2 ( .D(data[2]), .TD(q3_all[33]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[34]) );
  QDFZRBS fifo_mem_reg_5_1 ( .D(data[1]), .TD(q3_all[31]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[33]) );
  QDFZRBS fifo_mem_reg_4_31 ( .D(data[31]), .TD(q3_all[30]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[31]) );
  QDFZRBS fifo_mem_reg_4_28 ( .D(data[28]), .TD(q3_all[27]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[28]) );
  QDFZRBS fifo_mem_reg_4_27 ( .D(data[27]), .TD(q3_all[26]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[27]) );
  QDFZRBS fifo_mem_reg_4_26 ( .D(data[26]), .TD(q3_all[25]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[26]) );
  QDFZRBS fifo_mem_reg_4_25 ( .D(data[25]), .TD(q3_all[23]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[25]) );
  QDFZRBS fifo_mem_reg_4_23 ( .D(data[23]), .TD(q3_all[22]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[23]) );
  QDFZRBS fifo_mem_reg_4_22 ( .D(data[22]), .TD(q3_all[21]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[22]) );
  QDFZRBS fifo_mem_reg_4_19 ( .D(data[19]), .TD(q3_all[18]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[19]) );
  QDFZRBS fifo_mem_reg_4_18 ( .D(data[18]), .TD(q3_all[17]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[18]) );
  QDFZRBS fifo_mem_reg_4_17 ( .D(data[17]), .TD(q3_all[15]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[17]) );
  QDFZRBS fifo_mem_reg_4_15 ( .D(data[15]), .TD(q3_all[14]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[15]) );
  QDFZRBS fifo_mem_reg_4_14 ( .D(data[14]), .TD(q3_all[13]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[14]) );
  QDFZRBS fifo_mem_reg_4_11 ( .D(data[11]), .TD(q3_all[10]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[11]) );
  QDFZRBS fifo_mem_reg_4_10 ( .D(data[10]), .TD(q3_all[9]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[10]) );
  QDFZRBS fifo_mem_reg_4_9 ( .D(data[9]), .TD(q3_all[7]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[9])
         );
  QDFZRBS fifo_mem_reg_4_7 ( .D(data[7]), .TD(q3_all[6]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[7])
         );
  QDFZRBS fifo_mem_reg_4_6 ( .D(data[6]), .TD(q3_all[5]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[6])
         );
  QDFZRBS fifo_mem_reg_4_3 ( .D(data[3]), .TD(q3_all[2]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[3])
         );
  QDFZRBS fifo_mem_reg_4_2 ( .D(data[2]), .TD(q3_all[1]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[2])
         );
  QDFZRBS fifo_mem_reg_4_1 ( .D(data[1]), .TD(q2_all[63]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[1])
         );
  QDFZRBS fifo_mem_reg_1_30 ( .D(data[30]), .TD(q1_all[61]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[62]) );
  QDFZRBS fifo_mem_reg_1_29 ( .D(data[29]), .TD(q1_all[60]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[61]) );
  QDFZRBS fifo_mem_reg_1_14 ( .D(data[14]), .TD(q1_all[45]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N115_0_0), .RB(hresetn), .Q(
        q1_all[46]) );
  QDFZRBS fifo_mem_reg_0_30 ( .D(data[30]), .TD(q1_all[29]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[30]) );
  QDFZRBS fifo_mem_reg_0_21 ( .D(data[21]), .TD(q1_all[20]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[21]) );
  QDFZRBS fifo_mem_reg_0_13 ( .D(data[13]), .TD(q1_all[12]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[13]) );
  QDFZRBS fifo_mem_reg_0_12 ( .D(data[12]), .TD(q1_all[11]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(
        q1_all[12]) );
  QDFZRBS fifo_mem_reg_0_5 ( .D(data[5]), .TD(q1_all[4]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N83_0_0), .RB(hresetn), .Q(q1_all[5])
         );
  QDFZRBS fifo_mem_reg_5_30 ( .D(data[30]), .TD(q3_all[61]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[62]) );
  QDFZRBS fifo_mem_reg_5_29 ( .D(data[29]), .TD(q3_all[60]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[61]) );
  QDFZRBS fifo_mem_reg_5_22 ( .D(data[22]), .TD(q3_all[53]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[54]) );
  QDFZRBS fifo_mem_reg_5_14 ( .D(data[14]), .TD(q3_all[45]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[46]) );
  QDFZRBS fifo_mem_reg_5_13 ( .D(data[13]), .TD(q3_all[44]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(
        q3_all[45]) );
  QDFZRBS fifo_mem_reg_5_6 ( .D(data[6]), .TD(q3_all[37]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N243_0_0), .RB(hresetn), .Q(q3_all[38]) );
  QDFZRBS fifo_mem_reg_4_30 ( .D(data[30]), .TD(q3_all[29]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[30]) );
  QDFZRBS fifo_mem_reg_4_29 ( .D(data[29]), .TD(q3_all[28]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[29]) );
  QDFZRBS fifo_mem_reg_4_21 ( .D(data[21]), .TD(q3_all[20]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[21]) );
  QDFZRBS fifo_mem_reg_4_20 ( .D(data[20]), .TD(q3_all[19]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[20]) );
  QDFZRBS fifo_mem_reg_4_13 ( .D(data[13]), .TD(q3_all[12]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[13]) );
  QDFZRBS fifo_mem_reg_4_12 ( .D(data[12]), .TD(q3_all[11]), .SEL(test_se), 
        .CK(CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(
        q3_all[12]) );
  QDFZRBS fifo_mem_reg_4_5 ( .D(data[5]), .TD(q3_all[4]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[5])
         );
  QDFZRBS fifo_mem_reg_4_4 ( .D(data[4]), .TD(q3_all[3]), .SEL(test_se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N211_0_0), .RB(hresetn), .Q(q3_all[4])
         );
  QDFZRBS wr_ptr_reg_1 ( .D(n38), .TD(wr_ptr_0_), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(wr_ptr_1_) );
  QDFZRBS ptr_reg_1 ( .D(n41), .TD(ptr[0]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(ptr[1]) );
  QDFZRBS wr_ptr_reg_0 ( .D(n39), .TD(ptr[2]), .SEL(test_se), .CK(hclk), .RB(
        hresetn), .Q(wr_ptr_0_) );
  DFZRBS wr_ptr_reg_2 ( .D(n37), .TD(wr_ptr_1_), .SEL(test_se), .CK(hclk), 
        .RB(hresetn), .Q(test_so1), .QB(n11) );
  QDBHN LOCKUP ( .CKB(CLKGATING_hclk_POWERGATING_hclk_N147_0_0), .D(q2_all[15]), .Q(test_so2) );
endmodule


module des ( hclk, POR, hresetn, hsel, hwdata, haddr, hwrite, htrans, hsize, 
        hburst, hready, hready_resp, hresp, hrdata, Test_Mode, Test_Se, si0, 
        si1, si2, si3, so0, so1, so2, so3 );
  input [31:0] hwdata;
  input [9:0] haddr;
  input [1:0] htrans;
  input [2:0] hsize;
  input [2:0] hburst;
  output [1:0] hresp;
  output [31:0] hrdata;
  input hclk, POR, hresetn, hsel, hwrite, hready, Test_Mode, Test_Se, si0, si1,
         si2, si3;
  output hready_resp, so0, so1, so2, so3;
  wire   desctrl_sel, rw, desctrl_1, desctrl_0, run_delay, clr_ptr, desiv_sel,
         desiv_wr, deskey_sel, deskey_wr, desdat_rd, desdat_wr, des_start,
         desdat_full, nextiv_ready, nextiv_ready_en, desdat_ready, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, desctrl_sel_d1, desdat_sel_d1,
         deskey_sel_d1, desiv_sel_d1, N31, N32, N33, N34, N35, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N82, CLKGATING_hclk_POWERGATING_hclk_N26_0_0,
         net1749, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n24, n25, n26, n27, n29, n34, n35,
         n36, n37, n38, n39, n40, n41, n45, n48, n23, n31, n42, n43, n47, n49;
  wire   [31:0] dbusin;
  wire   [7:4] desctrl;
  wire   [1:0] edr;
  wire   [31:0] desdat_8_out;
  wire   [63:0] deskey1_64_out;
  wire   [63:0] deskey2_64_out;
  wire   [63:0] deskey3_64_out;
  wire   [63:0] desdat_64_out;
  wire   [63:0] desiv_64_out;
  wire   [63:0] desdat_64_in;

  NR2F U38 ( .I1(n7), .I2(n11), .O(n8) );
  des_key deskey_unit ( .hresetn(hresetn), .clrptr(clr_ptr), .hclk(hclk), .wr(
        deskey_wr), .data(dbusin), .q1_all(deskey1_64_out), .q2_all(
        deskey2_64_out), .q3_all(deskey3_64_out), .test_mode(Test_Mode), 
        .test_se(Test_Se), .test_si1(si3), .test_si2(deskey_sel), .test_so2(
        so2), .test_so1(n23) );
  des_iv desiv_unit ( .hclk(hclk), .POR(POR), .hresetn(hresetn), .clrptr(
        clr_ptr), .wr(desiv_wr), .deswr(nextiv_ready), .data(dbusin), 
        .data_all(desdat_64_out), .q_all(desiv_64_out), .test_mode(Test_Mode), 
        .test_se(Test_Se), .test_si1(si2), .test_si2(desiv_sel), .test_so2(so1), .test_so1(n31) );
  des_dat desdat_unit ( .POR(POR), .hresetn(hresetn), .clrptr(clr_ptr), .hclk(
        hclk), .rd(desdat_rd), .wr(desdat_wr), .deswr(desdat_ready), .data(
        dbusin), .data_all(desdat_64_in), .full_pulse(desdat_full), .q(
        desdat_8_out), .q_all(desdat_64_out), .test_mode(Test_Mode), .test_se(
        Test_Se), .test_si(n43), .test_so(n42) );
  des_cop des_cop_unit ( .hclk(hclk), .POR(POR), .hresetn(hresetn), 
        .encrypt_whole(desctrl[6]), .dt_sel(desctrl[5]), .key23_sel(desctrl[4]), .edr(edr), .mode_sel(desctrl_1), .iv_sel(desctrl_0), .iv(desiv_64_out), 
        .key1(deskey1_64_out), .key2(deskey2_64_out), .key3(deskey3_64_out), 
        .din(desdat_64_out), .din_valid_whole(des_start), .dout(desdat_64_in), 
        .dout_valid(desdat_ready), .test_mode(Test_Mode), .test_se(Test_Se), 
        .test_si(dbusin[31]), .test_so(n47) );
  POWERMODULE_HIGH_des_0 POWERGATING_hclk_N26_0 ( .CLK(hclk), .EN(N26), 
        .ENCLK(CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .TE(Test_Mode), 
        .ENOBS(net1749) );
  SNPS_CLOCK_GATE_OBS_des clk_gate_obs ( .TE(Test_Mode), .net1749(net1749), 
        .hclk(hclk), .test_se(Test_Se), .test_si(si0), .test_so(n49) );
  TIE1 U120 ( .O(n45) );
  INV2 U121 ( .I(n45), .O(hresp[0]) );
  INV2 U122 ( .I(n45), .O(hresp[1]) );
  ND2P U123 ( .I1(n11), .I2(n41), .O(n9) );
  NR2P U124 ( .I1(rw), .I2(n12), .O(desdat_wr) );
  ND3 U125 ( .I1(n4), .I2(n6), .I3(desctrl_sel), .O(n27) );
  OR3B2 U126 ( .I1(n48), .B1(n24), .B2(n25), .O(n5) );
  OR2 U127 ( .I1(haddr[6]), .I2(haddr[5]), .O(n48) );
  INV2 U128 ( .I(n13), .O(N32) );
  NR2 U129 ( .I1(n6), .I2(n12), .O(desdat_rd) );
  INV3 U130 ( .I(desdat_ready), .O(n4) );
  ND2 U131 ( .I1(n4), .I2(n27), .O(N26) );
  ND3P U132 ( .I1(n21), .I2(n22), .I3(n20), .O(n13) );
  OAI12S U133 ( .B1(n13), .B2(n16), .A1(n15), .O(N42) );
  OA12 U134 ( .B1(n13), .B2(n14), .A1(n15), .O(N82) );
  INV1 U135 ( .I(n18), .O(N34) );
  INV1 U136 ( .I(n19), .O(N33) );
  INV2 U137 ( .I(n17), .O(N35) );
  AOI112P U138 ( .C1(n5), .C2(n6), .A1(n7), .B1(N31), .O(n29) );
  NR2P U139 ( .I1(n14), .I2(n5), .O(N31) );
  INV2 U140 ( .I(n27), .O(n26) );
  AN2 U141 ( .I1(rw), .I2(desctrl_sel), .O(n11) );
  MOAI1 U142 ( .A1(n40), .A2(n9), .B1(desdat_8_out[0]), .B2(n8), .O(hrdata[0])
         );
  MOAI1 U143 ( .A1(n34), .A2(n9), .B1(desdat_8_out[1]), .B2(n8), .O(hrdata[1])
         );
  MOAI1 U144 ( .A1(n39), .A2(n9), .B1(desdat_8_out[2]), .B2(n8), .O(hrdata[2])
         );
  MOAI1 U145 ( .A1(n38), .A2(n9), .B1(desdat_8_out[3]), .B2(n8), .O(hrdata[3])
         );
  MOAI1 U146 ( .A1(n37), .A2(n9), .B1(desdat_8_out[4]), .B2(n8), .O(hrdata[4])
         );
  MOAI1 U147 ( .A1(n36), .A2(n9), .B1(desdat_8_out[5]), .B2(n8), .O(hrdata[5])
         );
  MOAI1 U148 ( .A1(n35), .A2(n9), .B1(desdat_8_out[6]), .B2(n8), .O(hrdata[6])
         );
  MOAI1 U149 ( .A1(n9), .A2(n10), .B1(desdat_8_out[7]), .B2(n8), .O(hrdata[7])
         );
  AN2 U150 ( .I1(desdat_8_out[10]), .I2(n8), .O(hrdata[10]) );
  AN2 U151 ( .I1(desdat_8_out[11]), .I2(n8), .O(hrdata[11]) );
  AN2 U152 ( .I1(desdat_8_out[12]), .I2(n8), .O(hrdata[12]) );
  AN2 U153 ( .I1(desdat_8_out[13]), .I2(n8), .O(hrdata[13]) );
  AN2 U154 ( .I1(desdat_8_out[14]), .I2(n8), .O(hrdata[14]) );
  AN2 U155 ( .I1(desdat_8_out[15]), .I2(n8), .O(hrdata[15]) );
  AN2 U156 ( .I1(desdat_8_out[16]), .I2(n8), .O(hrdata[16]) );
  AN2 U157 ( .I1(desdat_8_out[17]), .I2(n8), .O(hrdata[17]) );
  AN2 U158 ( .I1(desdat_8_out[18]), .I2(n8), .O(hrdata[18]) );
  AN2 U159 ( .I1(desdat_8_out[19]), .I2(n8), .O(hrdata[19]) );
  AN2 U160 ( .I1(desdat_8_out[20]), .I2(n8), .O(hrdata[20]) );
  AN2 U161 ( .I1(desdat_8_out[21]), .I2(n8), .O(hrdata[21]) );
  AN2 U162 ( .I1(desdat_8_out[22]), .I2(n8), .O(hrdata[22]) );
  AN2 U163 ( .I1(desdat_8_out[23]), .I2(n8), .O(hrdata[23]) );
  AN2 U164 ( .I1(desdat_8_out[24]), .I2(n8), .O(hrdata[24]) );
  AN2 U165 ( .I1(desdat_8_out[25]), .I2(n8), .O(hrdata[25]) );
  AN2 U166 ( .I1(desdat_8_out[26]), .I2(n8), .O(hrdata[26]) );
  AN2 U167 ( .I1(desdat_8_out[27]), .I2(n8), .O(hrdata[27]) );
  AN2 U168 ( .I1(desdat_8_out[28]), .I2(n8), .O(hrdata[28]) );
  AN2 U169 ( .I1(desdat_8_out[29]), .I2(n8), .O(hrdata[29]) );
  AN2 U170 ( .I1(desdat_8_out[30]), .I2(n8), .O(hrdata[30]) );
  AN2 U171 ( .I1(desdat_8_out[31]), .I2(n8), .O(hrdata[31]) );
  AN2 U172 ( .I1(desdat_8_out[8]), .I2(n8), .O(hrdata[8]) );
  AN2 U173 ( .I1(desdat_8_out[9]), .I2(n8), .O(hrdata[9]) );
  INV2 U174 ( .I(desctrl[7]), .O(n10) );
  AN2 U175 ( .I1(desiv_sel), .I2(n6), .O(desiv_wr) );
  NR2 U176 ( .I1(n3), .I2(n34), .O(nextiv_ready) );
  MAOI1 U177 ( .A1(nextiv_ready_en), .A2(n35), .B1(n35), .B2(n4), .O(n3) );
  AN2 U178 ( .I1(deskey_sel), .I2(n6), .O(deskey_wr) );
  NR3P U179 ( .I1(haddr[1]), .I2(haddr[0]), .I3(n5), .O(n20) );
  ND3 U180 ( .I1(n20), .I2(n21), .I3(haddr[3]), .O(n18) );
  ND3 U181 ( .I1(n20), .I2(n22), .I3(haddr[2]), .O(n19) );
  ND3 U182 ( .I1(haddr[2]), .I2(n20), .I3(haddr[3]), .O(n17) );
  AN4B1 U183 ( .I1(htrans[1]), .I2(hsel), .I3(hready), .B1(haddr[4]), .O(n25)
         );
  NR3P U184 ( .I1(haddr[7]), .I2(haddr[9]), .I3(haddr[8]), .O(n24) );
  MOAI1 U185 ( .A1(n16), .A2(n18), .B1(deskey_sel_d1), .B2(n7), .O(N44) );
  MOAI1 U186 ( .A1(n16), .A2(n19), .B1(desdat_sel_d1), .B2(n7), .O(N43) );
  MOAI1 U187 ( .A1(n16), .A2(n17), .B1(desiv_sel_d1), .B2(n7), .O(N45) );
  ND2P U188 ( .I1(n41), .I2(n14), .O(n16) );
  INV2 U189 ( .I(hwrite), .O(n14) );
  INV2 U190 ( .I(haddr[3]), .O(n22) );
  INV2 U191 ( .I(haddr[2]), .O(n21) );
  AN2 U192 ( .I1(hwdata[0]), .I2(n7), .O(N46) );
  AN2 U193 ( .I1(hwdata[1]), .I2(n7), .O(N47) );
  AN2 U194 ( .I1(hwdata[2]), .I2(n7), .O(N48) );
  AN2 U195 ( .I1(hwdata[3]), .I2(n7), .O(N49) );
  AN2 U196 ( .I1(hwdata[4]), .I2(n7), .O(N50) );
  AN2 U197 ( .I1(hwdata[5]), .I2(n7), .O(N51) );
  AN2 U198 ( .I1(hwdata[6]), .I2(n7), .O(N52) );
  AN2 U199 ( .I1(hwdata[7]), .I2(n7), .O(N53) );
  AN2 U200 ( .I1(hwdata[8]), .I2(n7), .O(N54) );
  AN2 U201 ( .I1(hwdata[9]), .I2(n7), .O(N55) );
  AN2 U202 ( .I1(hwdata[10]), .I2(n7), .O(N56) );
  AN2 U203 ( .I1(hwdata[11]), .I2(n7), .O(N57) );
  AN2 U204 ( .I1(hwdata[12]), .I2(n7), .O(N58) );
  AN2 U205 ( .I1(hwdata[13]), .I2(n7), .O(N59) );
  AN2 U206 ( .I1(hwdata[14]), .I2(n7), .O(N60) );
  AN2 U207 ( .I1(hwdata[15]), .I2(n7), .O(N61) );
  AN2 U208 ( .I1(hwdata[16]), .I2(n7), .O(N62) );
  AN2 U209 ( .I1(hwdata[17]), .I2(n7), .O(N63) );
  AN2 U210 ( .I1(hwdata[18]), .I2(n7), .O(N64) );
  AN2 U211 ( .I1(hwdata[19]), .I2(n7), .O(N65) );
  AN2 U212 ( .I1(hwdata[20]), .I2(n7), .O(N66) );
  AN2 U213 ( .I1(hwdata[21]), .I2(n7), .O(N67) );
  AN2 U214 ( .I1(hwdata[22]), .I2(n7), .O(N68) );
  AN2 U215 ( .I1(hwdata[23]), .I2(n7), .O(N69) );
  AN2 U216 ( .I1(hwdata[24]), .I2(n7), .O(N70) );
  AN2 U217 ( .I1(hwdata[25]), .I2(n7), .O(N71) );
  AN2 U218 ( .I1(hwdata[26]), .I2(n7), .O(N72) );
  AN2 U219 ( .I1(hwdata[27]), .I2(n7), .O(N73) );
  AN2 U220 ( .I1(hwdata[28]), .I2(n7), .O(N74) );
  AN2 U221 ( .I1(hwdata[29]), .I2(n7), .O(N75) );
  AN2 U222 ( .I1(hwdata[30]), .I2(n7), .O(N76) );
  AN2 U223 ( .I1(hwdata[31]), .I2(n7), .O(N77) );
  OR2P U224 ( .I1(run_delay), .I2(n10), .O(clr_ptr) );
  ND2 U225 ( .I1(desctrl_sel_d1), .I2(n7), .O(n15) );
  MOAI1 U226 ( .A1(n35), .A2(n4), .B1(dbusin[6]), .B2(n26), .O(N25) );
  MOAI1 U227 ( .A1(n34), .A2(n4), .B1(dbusin[1]), .B2(n26), .O(N20) );
  MOAI1 U228 ( .A1(n39), .A2(n4), .B1(dbusin[2]), .B2(n26), .O(N21) );
  MOAI1 U229 ( .A1(n38), .A2(n4), .B1(dbusin[3]), .B2(n26), .O(N22) );
  MOAI1 U230 ( .A1(n37), .A2(n4), .B1(dbusin[4]), .B2(n26), .O(N23) );
  MOAI1 U231 ( .A1(n36), .A2(n4), .B1(dbusin[5]), .B2(n26), .O(N24) );
  MOAI1 U232 ( .A1(n40), .A2(n4), .B1(dbusin[0]), .B2(n26), .O(N19) );
  AN2 U233 ( .I1(dbusin[7]), .I2(n26), .O(N27) );
  AN2 U234 ( .I1(desdat_full), .I2(desctrl[7]), .O(des_start) );
  des_spares_0 u_des_spares_0 ( .clk(hclk), .resetn(hresetn), .test_se(Test_Se), .test_si(rw), .test_so(so3) );
  QDFZRBS desdat_sel_d1_reg ( .D(N33), .TD(desctrl_sel), .SEL(Test_Se), .CK(
        hclk), .RB(hresetn), .Q(desdat_sel_d1) );
  QDFZRBS deskey_sel_d1_reg ( .D(N34), .TD(n31), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(deskey_sel_d1) );
  QDFZRBS desiv_sel_d1_reg ( .D(N35), .TD(n42), .SEL(Test_Se), .CK(hclk), .RB(
        hresetn), .Q(desiv_sel_d1) );
  QDFZRBS desctrl_sel_d1_reg ( .D(N32), .TD(desctrl[7]), .SEL(Test_Se), .CK(
        hclk), .RB(hresetn), .Q(desctrl_sel_d1) );
  QDFZRBS data_in_reg_24 ( .D(N70), .TD(dbusin[23]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[24]) );
  QDFZRBS data_in_reg_16 ( .D(N62), .TD(dbusin[15]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[16]) );
  QDFZRBS data_in_reg_8 ( .D(N54), .TD(dbusin[7]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[8]) );
  QDFZRBS data_in_reg_0 ( .D(N46), .TD(n49), .SEL(Test_Se), .CK(hclk), .RB(
        hresetn), .Q(dbusin[0]) );
  QDFZRBS data_in_reg_31 ( .D(N77), .TD(dbusin[30]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[31]) );
  QDFZRBS data_in_reg_30 ( .D(N76), .TD(dbusin[29]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[30]) );
  QDFZRBS data_in_reg_29 ( .D(N75), .TD(dbusin[28]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[29]) );
  QDFZRBS data_in_reg_28 ( .D(N74), .TD(dbusin[27]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[28]) );
  QDFZRBS data_in_reg_27 ( .D(N73), .TD(dbusin[26]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[27]) );
  QDFZRBS data_in_reg_26 ( .D(N72), .TD(dbusin[25]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[26]) );
  QDFZRBS data_in_reg_25 ( .D(N71), .TD(dbusin[24]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[25]) );
  QDFZRBS data_in_reg_23 ( .D(N69), .TD(dbusin[22]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[23]) );
  QDFZRBS data_in_reg_22 ( .D(N68), .TD(dbusin[21]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[22]) );
  QDFZRBS data_in_reg_21 ( .D(N67), .TD(dbusin[20]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[21]) );
  QDFZRBS data_in_reg_20 ( .D(N66), .TD(dbusin[19]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[20]) );
  QDFZRBS data_in_reg_19 ( .D(N65), .TD(dbusin[18]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[19]) );
  QDFZRBS data_in_reg_18 ( .D(N64), .TD(dbusin[17]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[18]) );
  QDFZRBS data_in_reg_17 ( .D(N63), .TD(dbusin[16]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[17]) );
  QDFZRBS data_in_reg_15 ( .D(N61), .TD(dbusin[14]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[15]) );
  QDFZRBS data_in_reg_14 ( .D(N60), .TD(dbusin[13]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[14]) );
  QDFZRBS data_in_reg_13 ( .D(N59), .TD(dbusin[12]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[13]) );
  QDFZRBS data_in_reg_12 ( .D(N58), .TD(dbusin[11]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[12]) );
  QDFZRBS data_in_reg_11 ( .D(N57), .TD(dbusin[10]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[11]) );
  QDFZRBS data_in_reg_10 ( .D(N56), .TD(dbusin[9]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[10]) );
  QDFZRBS data_in_reg_9 ( .D(N55), .TD(dbusin[8]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[9]) );
  QDFZRBS data_in_reg_7 ( .D(N53), .TD(dbusin[6]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[7]) );
  QDFZRBS data_in_reg_6 ( .D(N52), .TD(dbusin[5]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[6]) );
  QDFZRBS data_in_reg_5 ( .D(N51), .TD(dbusin[4]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[5]) );
  QDFZRBS data_in_reg_4 ( .D(N50), .TD(dbusin[3]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[4]) );
  QDFZRBS data_in_reg_3 ( .D(N49), .TD(dbusin[2]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[3]) );
  QDFZRBS data_in_reg_2 ( .D(N48), .TD(dbusin[1]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[2]) );
  QDFZRBS data_in_reg_1 ( .D(N47), .TD(dbusin[0]), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(dbusin[1]) );
  QDFZRBS run_delay_reg ( .D(desctrl[7]), .TD(nextiv_ready_en), .SEL(Test_Se), 
        .CK(hclk), .RB(hresetn), .Q(run_delay) );
  QDFZRBS deskey_sel_reg ( .D(N44), .TD(deskey_sel_d1), .SEL(Test_Se), .CK(
        hclk), .RB(hresetn), .Q(deskey_sel) );
  QDFZRBS nextiv_ready_en_reg ( .D(desdat_ready), .TD(n7), .SEL(Test_Se), .CK(
        hclk), .RB(hresetn), .Q(nextiv_ready_en) );
  QDFZRBS desiv_sel_reg ( .D(N45), .TD(desiv_sel_d1), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(desiv_sel) );
  QDFZRBS desctrl_reg_7 ( .D(N27), .TD(desctrl[6]), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(desctrl[7])
         );
  QDFZRBS desctrl_sel_reg ( .D(N42), .TD(desctrl_sel_d1), .SEL(Test_Se), .CK(
        hclk), .RB(hresetn), .Q(desctrl_sel) );
  DFZRBS desdat_sel_reg ( .D(N43), .TD(desdat_sel_d1), .SEL(Test_Se), .CK(hclk), .RB(hresetn), .Q(n43), .QB(n12) );
  DFZRBS desctrl_reg_6 ( .D(N25), .TD(desctrl[5]), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(desctrl[6]), 
        .QB(n35) );
  DFZRBS desctrl_reg_5 ( .D(N24), .TD(si1), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(desctrl[5]), 
        .QB(n36) );
  DFZRBS desctrl_reg_4 ( .D(N23), .TD(edr[1]), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(desctrl[4]), 
        .QB(n37) );
  DFZRBS desctrl_reg_3 ( .D(N22), .TD(edr[0]), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(edr[1]), 
        .QB(n38) );
  DFZRBS desctrl_reg_1 ( .D(N20), .TD(desctrl_0), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(desctrl_1), 
        .QB(n34) );
  DFZRBS desctrl_reg_0 ( .D(N19), .TD(n47), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(desctrl_0), 
        .QB(n40) );
  DFZRBS hwrite_d1_reg ( .D(N31), .TD(hready_resp), .SEL(Test_Se), .CK(hclk), 
        .RB(hresetn), .Q(n7), .QB(n41) );
  DFZSBN rw_reg ( .D(n29), .TD(run_delay), .SEL(Test_Se), .CK(hclk), .SB(
        hresetn), .Q(rw), .QB(n6) );
  DFZSBN hready_resp_reg ( .D(N82), .TD(n23), .SEL(Test_Se), .CK(hclk), .SB(
        hresetn), .Q(hready_resp) );
  DFZRBS desctrl_reg_2 ( .D(N21), .TD(desctrl_1), .SEL(Test_Se), .CK(
        CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .RB(hresetn), .Q(edr[0]), 
        .QB(n39) );
  QDBHN LOCKUP ( .CKB(CLKGATING_hclk_POWERGATING_hclk_N26_0_0), .D(desctrl[4]), 
        .Q(so0) );
endmodule

