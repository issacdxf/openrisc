// Verilog pattern output written by  TetraMAX (TM)  Z-2007.03-SP1-i070413_172030 
// Date: Fri Sep 18 17:15:31 2009
// Module tested: des

//     Uncollapsed Stuck Fault Summary Report
// -----------------------------------------------
// fault class                     code   #faults
// ------------------------------  ----  ---------
// Detected                         DT      34438
// Possibly detected                PT          0
// Undetectable                     UD        111
// ATPG untestable                  AU        546
// Not detected                     ND         13
// -----------------------------------------------
// total faults                             35108
// test coverage                            98.40%
// -----------------------------------------------
// 
//            Pattern Summary Report
// -----------------------------------------------
// #internal patterns                         131
//     #basic_scan patterns                   131
// -----------------------------------------------
// 
// rule  severity  #fails  description
// ----  --------  ------  ---------------------------------
// N2    warning      128  unsupported construct
// N16   warning        1  overspecified UDP
// N23   warning        1  inconsistent UDP
// B8    warning       20  unconnected module input pin
// B9    warning        1  undriven module internal net
// B10   warning        4  unconnected module internal net
// 
// clock_name        off  usage
// ----------------  ---  --------------------------
// hclk               0   master shift nonscan_DLAT 
// 
// port_name         constraint_value
// ----------------  ---------------
// POR                 1
// hresetn             1
// Test_Mode           1
// 
// There are no equivalent pins
// There are no net connections

`timescale 1 ns / 1 ns

//
// --- NOTE: Remove the comment to define 'tmax_iddq' to activate processing of IDDQ events
//     Or use '+define+tmax_iddq' on the verilog compile line
//
//`define tmax_iddq

module AAA_tmax_testbench_1_16 ;
   parameter NAMELENGTH = 200; // max length of names reported in fails
   parameter LENMAX = 112, NSHIFTS = 1; // LENMAX for serial
   parameter LENSERIAL = 112, NCHAINS = 4;
   parameter SHBEG = 0, SHEND = 0;
   integer nofails, bit, cbit, pattern, lastpattern, chain, idx;
   integer error_banner; // flag for tracking displayed error banner
   integer loads;        // number of load_unloads for current pattern
   integer patm1;        // pattern - 1
   integer patp1;        // pattern + lastpattern
   integer prev_pat;     // previous pattern number
   integer report_interval; // report pattern progress every Nth pattern
   integer verbose;      // message verbosity level
   parameter NINPUTS = 62, NOUTPUTS = 39;
   wire [0:NOUTPUTS-1] PO; reg [0:NOUTPUTS-1] ALLPOS, XPCT, MASK;
   reg [0:NINPUTS-1] PI, ALLPIS;
   reg [0:8*(NAMELENGTH-1)] POnames [0:NOUTPUTS-1];
   reg [0:8*(NAMELENGTH-1)] CHAINnames [0:NCHAINS-1];
   reg [0:8*(NAMELENGTH-1)] CHAINpins [0:NCHAINS-1];
   reg [0:LENSERIAL-1] LOAD0, LOADSH0, LOAD1, LOADSH1, LOAD2, LOADSH2, LOAD3,
   LOADSH3;
   reg [0:LENMAX-1] UNL, UNLOAD[0:NCHAINS-1];
   reg [0:LENMAX-1] UNLM, UNLMSK[0:NCHAINS-1], SHBEGM[0:NCHAINS-1];
   reg [0:LENMAX-1] SERIALM;
   reg [0:LENMAX-1] INPINV[0:NCHAINS-1], OUTINV[0:NCHAINS-1];
   wire [0:NCHAINS-1] SCANOUT;
   wire [0:LENMAX-1] CHAINOUT0, CHAINOUT1, CHAINOUT2, CHAINOUT3;
   reg [0:LENMAX-1] CHOUT, CHAINOUT[0:NCHAINS-1];
   event IDDQ;

   wire hclk;
   wire POR;
   wire hresetn;
   wire hsel;
   wire hwrite;
   wire hready;
   wire hready_resp;
   wire Test_Mode;
   wire Test_Se;
   wire si0;
   wire si1;
   wire si2;
   wire si3;
   wire so0;
   wire so1;
   wire so2;
   wire so3;
   wire [31:0] hwdata;
   wire [9:0] haddr;
   wire [1:0] htrans;
   wire [2:0] hsize;
   wire [2:0] hburst;
   wire [1:0] hresp;
   wire [31:0] hrdata;

   // map PI[] vector to DUT inputs and bidis
   assign hclk = PI[0];
   assign POR = PI[1];
   assign hresetn = PI[2];
   assign hsel = PI[3];
   assign hwdata = PI[4:35];
   assign haddr = PI[36:45];
   assign hwrite = PI[46];
   assign htrans = PI[47:48];
   assign hsize = PI[49:51];
   assign hburst = PI[52:54];
   assign hready = PI[55];
   assign Test_Mode = PI[56];
   assign Test_Se = PI[57];
   assign si0 = PI[58];
   assign si1 = PI[59];
   assign si2 = PI[60];
   assign si3 = PI[61];

   // map DUT outputs and bidis to PO[] vector
   assign
      PO[0] = hready_resp ,
      PO[1] = hresp[1] ,
      PO[2] = hresp[0] ,
      PO[3] = hrdata[31] ,
      PO[4] = hrdata[30] ,
      PO[5] = hrdata[29] ,
      PO[6] = hrdata[28] ,
      PO[7] = hrdata[27] ,
      PO[8] = hrdata[26] ,
      PO[9] = hrdata[25] ,
      PO[10] = hrdata[24] ,
      PO[11] = hrdata[23] ,
      PO[12] = hrdata[22] ,
      PO[13] = hrdata[21] ,
      PO[14] = hrdata[20] ,
      PO[15] = hrdata[19] ,
      PO[16] = hrdata[18] ,
      PO[17] = hrdata[17] ,
      PO[18] = hrdata[16] ,
      PO[19] = hrdata[15] ,
      PO[20] = hrdata[14] ,
      PO[21] = hrdata[13] ,
      PO[22] = hrdata[12] ,
      PO[23] = hrdata[11] ,
      PO[24] = hrdata[10] ,
      PO[25] = hrdata[9] ,
      PO[26] = hrdata[8] ,
      PO[27] = hrdata[7] ,
      PO[28] = hrdata[6] ,
      PO[29] = hrdata[5] ,
      PO[30] = hrdata[4] ,
      PO[31] = hrdata[3] ;
   assign
      PO[32] = hrdata[2] ,
      PO[33] = hrdata[1] ,
      PO[34] = hrdata[0] ,
      PO[35] = so0 ,
      PO[36] = so1 ,
      PO[37] = so2 ,
      PO[38] = so3 ;

   // instantiate the design into the testbench
   des dut (
      .hclk(hclk),
      .POR(POR),
      .hresetn(hresetn),
      .hsel(hsel),
      .hwdata(hwdata),
      .haddr(haddr),
      .hwrite(hwrite),
      .htrans(htrans),
      .hsize(hsize),
      .hburst(hburst),
      .hready(hready),
      .hready_resp(hready_resp),
      .hresp(hresp),
      .hrdata(hrdata),
      .Test_Mode(Test_Mode),
      .Test_Se(Test_Se),
      .si0(si0),
      .si1(si1),
      .si2(si2),
      .si3(si3),
      .so0(so0),
      .so1(so1),
      .so2(so2),
      .so3(so3)   );

   event pulse_hclk;
   always @ pulse_hclk begin
      #45 PI[0] = 1; #10 PI[0] = 0;   // hclk
   end


   integer errshown;
   event measurePO;
   always @ measurePO begin
      if (((XPCT&MASK) !== (ALLPOS&MASK)) || (XPCT !== (~(~XPCT)))) begin
         errshown = 0;
         for (bit = 0; bit < NOUTPUTS; bit=bit + 1) begin
            if (MASK[bit]==1'b1) begin
               if (XPCT[bit] !== ALLPOS[bit]) begin
                  if (errshown==0) $display("\n// *** ERROR during capture pattern %0d, T=%t", pattern, $time);
                  $display("  %0d %0s (exp=%b, got=%b)", pattern, POnames[bit], XPCT[bit], ALLPOS[bit]);
                  nofails = nofails + 1; errshown = 1;
               end
            end
         end
      end
   end

   event forcePI_default_WFT;
   always @ forcePI_default_WFT begin
      PI = ALLPIS;
   end
   event measurePO_default_WFT;
   always @ measurePO_default_WFT begin
      #40;
      ALLPOS = PO;
      #0; #0 -> measurePO;
      `ifdef tmax_iddq
         #0; ->IDDQ;
      `endif
   end

   event force_scanin;
   always @ force_scanin begin
      PI[58] <= LOAD0[bit];
      PI[59] <= LOAD1[bit];
      PI[60] <= LOAD2[bit];
      PI[61] <= LOAD3[bit];
   end

   assign SCANOUT[0] = so0,  SCANOUT[1] = so1,  SCANOUT[2] = so2,  SCANOUT[3] = so3;

   event measure_scanout;
   always @ measure_scanout begin
      if ((NSHIFTS < LENMAX) && (bit >= SHBEG)) cbit = bit - LENMAX + NSHIFTS + 1 + SHBEG;
      else cbit = bit; // because parallel does NSHIFTS + 1 shifts
      idx = cbit + 0;
      for (chain = 0; chain < 4; chain=chain + 1) begin
         UNL = UNLOAD[chain]; UNLM = UNLMSK[chain];
         if ((UNL[idx]&UNLM[idx]) !== (SCANOUT[chain]&UNLM[idx])) begin
            patp1 = pattern + lastpattern;  patm1 = patp1 - 1;
            if (error_banner != pattern) begin
               if (lastpattern == 0) $display("\n// *** ERROR during scan pattern %0d (detected during load of pattern %0d)", patm1, patp1);
               else $display("\n// *** ERROR during scan pattern %0d (detected during final pattern unload)", patm1);
               error_banner = pattern;
            end
            $display("  %0d %0s %0d (exp=%b, got=%b)  // pin %0s, scan cell %0d, T=%t",
               patm1, CHAINnames[chain], cbit, UNL[idx], SCANOUT[chain], CHAINpins[chain], cbit, $time);
            nofails = nofails + 1;
         end
      end
   end


   always @ IDDQ begin
   `ifdef tmax_iddq
      $ssi_iddq("strobe_try");
      $ssi_iddq("status drivers leaky AAA_tmax_testbench_1_16.leaky");
   `endif
   end

   event capture;
   always @ capture begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
   end

   event capture_hclk;
   always @ capture_hclk begin
      ->forcePI_default_WFT;
      #100; ->measurePO_default_WFT;
      #145 PI[0] = 1; // hclk
      #10 PI[0] = 0; // hclk
   end

   task shift;
   begin
      if (verbose >= 4) $display("// %t :    shift %0d", $time, bit);
      ->force_scanin;
      #40; ->measure_scanout;
      #5 PI[0] = 1; // hclk
      #10 PI[0] = 0; // hclk
      #45;
   end
   endtask

   event test_setup;
   always @ test_setup begin
      #0 PI[1] = 1; // POR
      #0 PI[56] = 1; // Test_Mode
      #0 PI[0] = 0; // hclk
      #0 PI[2] = 1; // hresetn
      #0 PI[45] = 1'bX; // haddr[0]
      #0 PI[44] = 1'bX; // haddr[1]
      #0 PI[43] = 1'bX; // haddr[2]
      #0 PI[42] = 1'bX; // haddr[3]
      #0 PI[41] = 1'bX; // haddr[4]
      #0 PI[40] = 1'bX; // haddr[5]
      #0 PI[39] = 1'bX; // haddr[6]
      #0 PI[38] = 1'bX; // haddr[7]
      #0 PI[37] = 1'bX; // haddr[8]
      #0 PI[36] = 1'bX; // haddr[9]
      #0 PI[54] = 1'bX; // hburst[0]
      #0 PI[53] = 1'bX; // hburst[1]
      #0 PI[52] = 1'bX; // hburst[2]
      #0 PI[55] = 1'bX; // hready
      #0 PI[3] = 1'bX; // hsel
      #0 PI[51] = 1'bX; // hsize[0]
      #0 PI[50] = 1'bX; // hsize[1]
      #0 PI[49] = 1'bX; // hsize[2]
      #0 PI[48] = 1'bX; // htrans[0]
      #0 PI[47] = 1'bX; // htrans[1]
      #0 PI[35] = 1'bX; // hwdata[0]
      #0 PI[25] = 1'bX; // hwdata[10]
      #0 PI[24] = 1'bX; // hwdata[11]
      #0 PI[23] = 1'bX; // hwdata[12]
      #0 PI[22] = 1'bX; // hwdata[13]
      #0 PI[21] = 1'bX; // hwdata[14]
      #0 PI[20] = 1'bX; // hwdata[15]
      #0 PI[19] = 1'bX; // hwdata[16]
      #0 PI[18] = 1'bX; // hwdata[17]
      #0 PI[17] = 1'bX; // hwdata[18]
      #0 PI[16] = 1'bX; // hwdata[19]
      #0 PI[34] = 1'bX; // hwdata[1]
      #0 PI[15] = 1'bX; // hwdata[20]
      #0 PI[14] = 1'bX; // hwdata[21]
      #0 PI[13] = 1'bX; // hwdata[22]
      #0 PI[12] = 1'bX; // hwdata[23]
      #0 PI[11] = 1'bX; // hwdata[24]
      #0 PI[10] = 1'bX; // hwdata[25]
      #0 PI[9] = 1'bX; // hwdata[26]
      #0 PI[8] = 1'bX; // hwdata[27]
      #0 PI[7] = 1'bX; // hwdata[28]
      #0 PI[6] = 1'bX; // hwdata[29]
      #0 PI[33] = 1'bX; // hwdata[2]
      #0 PI[5] = 1'bX; // hwdata[30]
      #0 PI[4] = 1'bX; // hwdata[31]
      #0 PI[32] = 1'bX; // hwdata[3]
      #0 PI[31] = 1'bX; // hwdata[4]
      #0 PI[30] = 1'bX; // hwdata[5]
      #0 PI[29] = 1'bX; // hwdata[6]
      #0 PI[28] = 1'bX; // hwdata[7]
      #0 PI[27] = 1'bX; // hwdata[8]
      #0 PI[26] = 1'bX; // hwdata[9]
      #0 PI[46] = 1'bX; // hwrite
      #0 PI[57] = 1'bX; // Test_Se
      #0 PI[58] = 1'bX; // si0
      #0 PI[59] = 1'bX; // si1
      #0 PI[60] = 1'bX; // si2
      #0 PI[61] = 1'bX; // si3
   end


   task multiple_shift;
   begin
      bit = bit-1;
      error_banner = -2;
      while (bit+1 < LENMAX-SHEND) begin
         bit = bit+1;
         shift;
      end
   end
   endtask

   assign CHAINOUT0 = { dut.LOCKUP.Q, dut.desctrl_reg_3.Q, dut.desctrl_reg_2.Q, dut.desctrl_reg_1.Q,
          dut.desctrl_reg_0.Q, dut.des_cop_unit.flag_reg_1.Q, dut.des_cop_unit.flag_reg_0.Q,
          dut.des_cop_unit.din_valid_eins_reg.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_63.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_62.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_61.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_60.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_59.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_58.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_57.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_56.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_55.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_54.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_53.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_52.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_51.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_50.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_49.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_48.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_47.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_46.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_45.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_44.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_43.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_42.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_41.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_40.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_39.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_38.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_37.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_36.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_35.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_34.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_33.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_32.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_31.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_30.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_29.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_28.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_27.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_26.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_25.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_24.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_23.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_22.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_21.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_20.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_19.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_18.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_17.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_16.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_15.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_14.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_13.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_12.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_11.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_10.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_9.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_8.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_7.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_6.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_5.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_4.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_3.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_2.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_1.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_0.Q, 
          dut.des_cop_unit.des_unit.u_tiny_des_round.clk_gate_obs.U1.Q, 
          dut.des_cop_unit.des_unit.state_reg.Q, dut.des_cop_unit.des_unit.round_reg_3.Q,
          dut.des_cop_unit.des_unit.round_reg_2.Q, dut.des_cop_unit.des_unit.round_reg_1.Q,
          dut.des_cop_unit.des_unit.round_reg_0.Q, dut.des_cop_unit.des_unit.dout_valid_reg.Q,
          dut.data_in_reg_31.Q, dut.data_in_reg_30.Q, dut.data_in_reg_29.Q, dut.data_in_reg_28.Q,
          dut.data_in_reg_27.Q, dut.data_in_reg_26.Q, dut.data_in_reg_25.Q, dut.data_in_reg_24.Q,
          dut.data_in_reg_23.Q, dut.data_in_reg_22.Q, dut.data_in_reg_21.Q, dut.data_in_reg_20.Q,
          dut.data_in_reg_19.Q, dut.data_in_reg_18.Q, dut.data_in_reg_17.Q, dut.data_in_reg_16.Q,
          dut.data_in_reg_15.Q, dut.data_in_reg_14.Q, dut.data_in_reg_13.Q, dut.data_in_reg_12.Q,
          dut.data_in_reg_11.Q, dut.data_in_reg_10.Q, dut.data_in_reg_9.Q, dut.data_in_reg_8.Q,
          dut.data_in_reg_7.Q, dut.data_in_reg_6.Q, dut.data_in_reg_5.Q, dut.data_in_reg_4.Q,
          dut.data_in_reg_3.Q, dut.data_in_reg_2.Q, dut.data_in_reg_1.Q, dut.data_in_reg_0.Q,
          dut.clk_gate_obs.U1.Q };
   assign CHAINOUT1 = { dut.desiv_unit.LOCKUP.Q, dut.desiv_unit.fifo_mem_reg_0_27.Q,
          dut.desiv_unit.fifo_mem_reg_0_26.Q, dut.desiv_unit.fifo_mem_reg_0_25.Q,
          dut.desiv_unit.fifo_mem_reg_0_24.Q, dut.desiv_unit.fifo_mem_reg_0_23.Q,
          dut.desiv_unit.fifo_mem_reg_0_22.Q, dut.desiv_unit.fifo_mem_reg_0_21.Q,
          dut.desiv_unit.fifo_mem_reg_0_20.Q, dut.desiv_unit.fifo_mem_reg_0_19.Q,
          dut.desiv_unit.fifo_mem_reg_0_18.Q, dut.desiv_unit.fifo_mem_reg_0_17.Q,
          dut.desiv_unit.fifo_mem_reg_0_16.Q, dut.desiv_unit.fifo_mem_reg_0_15.Q,
          dut.desiv_unit.fifo_mem_reg_0_14.Q, dut.desiv_unit.fifo_mem_reg_0_13.Q,
          dut.desiv_unit.fifo_mem_reg_0_12.Q, dut.desiv_unit.fifo_mem_reg_0_11.Q,
          dut.desiv_unit.fifo_mem_reg_0_10.Q, dut.desiv_unit.fifo_mem_reg_0_9.Q,
          dut.desiv_unit.fifo_mem_reg_0_8.Q, dut.desiv_unit.fifo_mem_reg_0_7.Q, 
          dut.desiv_unit.fifo_mem_reg_0_6.Q, dut.desiv_unit.fifo_mem_reg_0_5.Q, 
          dut.desiv_unit.fifo_mem_reg_0_4.Q, dut.desiv_unit.fifo_mem_reg_0_3.Q, 
          dut.desiv_unit.fifo_mem_reg_0_2.Q, dut.desiv_unit.fifo_mem_reg_0_1.Q, 
          dut.desiv_unit.fifo_mem_reg_0_0.Q, dut.desiv_unit.clk_gate_obs.U1.Q, dut.desiv_sel_reg.Q,
          dut.desiv_sel_d1_reg.Q, dut.desdat_unit.wr_ptr_reg.Q, dut.desdat_unit.rd_ptr_reg.Q,
          dut.desdat_unit.ptr_reg_1.Q, dut.desdat_unit.ptr_reg_0.Q, dut.desdat_unit.full_reg.Q,
          dut.desdat_unit.full_pulse_reg.Q, dut.desdat_unit.full_delay_reg.Q, 
          dut.desdat_unit.fifo_mem_reg_1_31.Q, dut.desdat_unit.fifo_mem_reg_1_30.Q,
          dut.desdat_unit.fifo_mem_reg_1_29.Q, dut.desdat_unit.fifo_mem_reg_1_28.Q,
          dut.desdat_unit.fifo_mem_reg_1_27.Q, dut.desdat_unit.fifo_mem_reg_1_26.Q,
          dut.desdat_unit.fifo_mem_reg_1_25.Q, dut.desdat_unit.fifo_mem_reg_1_24.Q,
          dut.desdat_unit.fifo_mem_reg_1_23.Q, dut.desdat_unit.fifo_mem_reg_1_22.Q,
          dut.desdat_unit.fifo_mem_reg_1_21.Q, dut.desdat_unit.fifo_mem_reg_1_20.Q,
          dut.desdat_unit.fifo_mem_reg_1_19.Q, dut.desdat_unit.fifo_mem_reg_1_18.Q,
          dut.desdat_unit.fifo_mem_reg_1_17.Q, dut.desdat_unit.fifo_mem_reg_1_16.Q,
          dut.desdat_unit.fifo_mem_reg_1_15.Q, dut.desdat_unit.fifo_mem_reg_1_14.Q,
          dut.desdat_unit.fifo_mem_reg_1_13.Q, dut.desdat_unit.fifo_mem_reg_1_12.Q,
          dut.desdat_unit.fifo_mem_reg_1_11.Q, dut.desdat_unit.fifo_mem_reg_1_10.Q,
          dut.desdat_unit.fifo_mem_reg_1_9.Q, dut.desdat_unit.fifo_mem_reg_1_8.Q,
          dut.desdat_unit.fifo_mem_reg_1_7.Q, dut.desdat_unit.fifo_mem_reg_1_6.Q,
          dut.desdat_unit.fifo_mem_reg_1_5.Q, dut.desdat_unit.fifo_mem_reg_1_4.Q,
          dut.desdat_unit.fifo_mem_reg_1_3.Q, dut.desdat_unit.fifo_mem_reg_1_2.Q,
          dut.desdat_unit.fifo_mem_reg_1_1.Q, dut.desdat_unit.fifo_mem_reg_1_0.Q,
          dut.desdat_unit.fifo_mem_reg_0_31.Q, dut.desdat_unit.fifo_mem_reg_0_30.Q,
          dut.desdat_unit.fifo_mem_reg_0_29.Q, dut.desdat_unit.fifo_mem_reg_0_28.Q,
          dut.desdat_unit.fifo_mem_reg_0_27.Q, dut.desdat_unit.fifo_mem_reg_0_26.Q,
          dut.desdat_unit.fifo_mem_reg_0_25.Q, dut.desdat_unit.fifo_mem_reg_0_24.Q,
          dut.desdat_unit.fifo_mem_reg_0_23.Q, dut.desdat_unit.fifo_mem_reg_0_22.Q,
          dut.desdat_unit.fifo_mem_reg_0_21.Q, dut.desdat_unit.fifo_mem_reg_0_20.Q,
          dut.desdat_unit.fifo_mem_reg_0_19.Q, dut.desdat_unit.fifo_mem_reg_0_18.Q,
          dut.desdat_unit.fifo_mem_reg_0_17.Q, dut.desdat_unit.fifo_mem_reg_0_16.Q,
          dut.desdat_unit.fifo_mem_reg_0_15.Q, dut.desdat_unit.fifo_mem_reg_0_14.Q,
          dut.desdat_unit.fifo_mem_reg_0_13.Q, dut.desdat_unit.fifo_mem_reg_0_12.Q,
          dut.desdat_unit.fifo_mem_reg_0_11.Q, dut.desdat_unit.fifo_mem_reg_0_10.Q,
          dut.desdat_unit.fifo_mem_reg_0_9.Q, dut.desdat_unit.fifo_mem_reg_0_8.Q,
          dut.desdat_unit.fifo_mem_reg_0_7.Q, dut.desdat_unit.fifo_mem_reg_0_6.Q,
          dut.desdat_unit.fifo_mem_reg_0_5.Q, dut.desdat_unit.fifo_mem_reg_0_4.Q,
          dut.desdat_unit.fifo_mem_reg_0_3.Q, dut.desdat_unit.fifo_mem_reg_0_2.Q,
          dut.desdat_unit.fifo_mem_reg_0_1.Q, dut.desdat_unit.fifo_mem_reg_0_0.Q,
          dut.desdat_unit.clk_gate_obs.U1.Q, dut.desdat_sel_reg.Q, dut.desdat_sel_d1_reg.Q,
          dut.desctrl_sel_reg.Q, dut.desctrl_sel_d1_reg.Q, dut.desctrl_reg_7.Q, dut.desctrl_reg_6.Q,
          dut.desctrl_reg_5.Q, 1'b0 };
   assign CHAINOUT2 = { dut.deskey_unit.LOCKUP.Q, dut.deskey_unit.fifo_mem_reg_2_14.Q,
          dut.deskey_unit.fifo_mem_reg_2_13.Q, dut.deskey_unit.fifo_mem_reg_2_12.Q,
          dut.deskey_unit.fifo_mem_reg_2_11.Q, dut.deskey_unit.fifo_mem_reg_2_10.Q,
          dut.deskey_unit.fifo_mem_reg_2_9.Q, dut.deskey_unit.fifo_mem_reg_2_7.Q,
          dut.deskey_unit.fifo_mem_reg_2_6.Q, dut.deskey_unit.fifo_mem_reg_2_5.Q,
          dut.deskey_unit.fifo_mem_reg_2_4.Q, dut.deskey_unit.fifo_mem_reg_2_3.Q,
          dut.deskey_unit.fifo_mem_reg_2_2.Q, dut.deskey_unit.fifo_mem_reg_2_1.Q,
          dut.deskey_unit.fifo_mem_reg_1_31.Q, dut.deskey_unit.fifo_mem_reg_1_30.Q,
          dut.deskey_unit.fifo_mem_reg_1_29.Q, dut.deskey_unit.fifo_mem_reg_1_28.Q,
          dut.deskey_unit.fifo_mem_reg_1_27.Q, dut.deskey_unit.fifo_mem_reg_1_26.Q,
          dut.deskey_unit.fifo_mem_reg_1_25.Q, dut.deskey_unit.fifo_mem_reg_1_23.Q,
          dut.deskey_unit.fifo_mem_reg_1_22.Q, dut.deskey_unit.fifo_mem_reg_1_21.Q,
          dut.deskey_unit.fifo_mem_reg_1_20.Q, dut.deskey_unit.fifo_mem_reg_1_19.Q,
          dut.deskey_unit.fifo_mem_reg_1_18.Q, dut.deskey_unit.fifo_mem_reg_1_17.Q,
          dut.deskey_unit.fifo_mem_reg_1_15.Q, dut.deskey_unit.fifo_mem_reg_1_14.Q,
          dut.deskey_unit.fifo_mem_reg_1_13.Q, dut.deskey_unit.fifo_mem_reg_1_12.Q,
          dut.deskey_unit.fifo_mem_reg_1_11.Q, dut.deskey_unit.fifo_mem_reg_1_10.Q,
          dut.deskey_unit.fifo_mem_reg_1_9.Q, dut.deskey_unit.fifo_mem_reg_1_7.Q,
          dut.deskey_unit.fifo_mem_reg_1_6.Q, dut.deskey_unit.fifo_mem_reg_1_5.Q,
          dut.deskey_unit.fifo_mem_reg_1_4.Q, dut.deskey_unit.fifo_mem_reg_1_3.Q,
          dut.deskey_unit.fifo_mem_reg_1_2.Q, dut.deskey_unit.fifo_mem_reg_1_1.Q,
          dut.deskey_unit.fifo_mem_reg_0_31.Q, dut.deskey_unit.fifo_mem_reg_0_30.Q,
          dut.deskey_unit.fifo_mem_reg_0_29.Q, dut.deskey_unit.fifo_mem_reg_0_28.Q,
          dut.deskey_unit.fifo_mem_reg_0_27.Q, dut.deskey_unit.fifo_mem_reg_0_26.Q,
          dut.deskey_unit.fifo_mem_reg_0_25.Q, dut.deskey_unit.fifo_mem_reg_0_23.Q,
          dut.deskey_unit.fifo_mem_reg_0_22.Q, dut.deskey_unit.fifo_mem_reg_0_21.Q,
          dut.deskey_unit.fifo_mem_reg_0_20.Q, dut.deskey_unit.fifo_mem_reg_0_19.Q,
          dut.deskey_unit.fifo_mem_reg_0_18.Q, dut.deskey_unit.fifo_mem_reg_0_17.Q,
          dut.deskey_unit.fifo_mem_reg_0_15.Q, dut.deskey_unit.fifo_mem_reg_0_14.Q,
          dut.deskey_unit.fifo_mem_reg_0_13.Q, dut.deskey_unit.fifo_mem_reg_0_12.Q,
          dut.deskey_unit.fifo_mem_reg_0_11.Q, dut.deskey_unit.fifo_mem_reg_0_10.Q,
          dut.deskey_unit.fifo_mem_reg_0_9.Q, dut.deskey_unit.fifo_mem_reg_0_7.Q,
          dut.deskey_unit.fifo_mem_reg_0_6.Q, dut.deskey_unit.fifo_mem_reg_0_5.Q,
          dut.deskey_unit.fifo_mem_reg_0_4.Q, dut.deskey_unit.fifo_mem_reg_0_3.Q,
          dut.deskey_unit.fifo_mem_reg_0_2.Q, dut.deskey_unit.fifo_mem_reg_0_1.Q,
          dut.deskey_unit.clk_gate_obs.U1.Q, dut.deskey_sel_reg.Q, dut.deskey_sel_d1_reg.Q,
          dut.desiv_unit.wr_ptr_reg.Q, dut.desiv_unit.ptr_reg_1.Q, dut.desiv_unit.ptr_reg_0.Q,
          dut.desiv_unit.fifo_mem_reg_1_31.Q, dut.desiv_unit.fifo_mem_reg_1_30.Q,
          dut.desiv_unit.fifo_mem_reg_1_29.Q, dut.desiv_unit.fifo_mem_reg_1_28.Q,
          dut.desiv_unit.fifo_mem_reg_1_27.Q, dut.desiv_unit.fifo_mem_reg_1_26.Q,
          dut.desiv_unit.fifo_mem_reg_1_25.Q, dut.desiv_unit.fifo_mem_reg_1_24.Q,
          dut.desiv_unit.fifo_mem_reg_1_23.Q, dut.desiv_unit.fifo_mem_reg_1_22.Q,
          dut.desiv_unit.fifo_mem_reg_1_21.Q, dut.desiv_unit.fifo_mem_reg_1_20.Q,
          dut.desiv_unit.fifo_mem_reg_1_19.Q, dut.desiv_unit.fifo_mem_reg_1_18.Q,
          dut.desiv_unit.fifo_mem_reg_1_17.Q, dut.desiv_unit.fifo_mem_reg_1_16.Q,
          dut.desiv_unit.fifo_mem_reg_1_15.Q, dut.desiv_unit.fifo_mem_reg_1_14.Q,
          dut.desiv_unit.fifo_mem_reg_1_13.Q, dut.desiv_unit.fifo_mem_reg_1_12.Q,
          dut.desiv_unit.fifo_mem_reg_1_11.Q, dut.desiv_unit.fifo_mem_reg_1_10.Q,
          dut.desiv_unit.fifo_mem_reg_1_9.Q, dut.desiv_unit.fifo_mem_reg_1_8.Q, 
          dut.desiv_unit.fifo_mem_reg_1_7.Q, dut.desiv_unit.fifo_mem_reg_1_6.Q, 
          dut.desiv_unit.fifo_mem_reg_1_5.Q, dut.desiv_unit.fifo_mem_reg_1_4.Q, 
          dut.desiv_unit.fifo_mem_reg_1_3.Q, dut.desiv_unit.fifo_mem_reg_1_2.Q, 
          dut.desiv_unit.fifo_mem_reg_1_1.Q, dut.desiv_unit.fifo_mem_reg_1_0.Q, 
          dut.desiv_unit.fifo_mem_reg_0_31.Q, dut.desiv_unit.fifo_mem_reg_0_30.Q,
          dut.desiv_unit.fifo_mem_reg_0_29.Q, 1'b0 };
   assign CHAINOUT3 = { dut.u_des_spares_0.LOCKUP.Q, dut.u_des_spares_0.SPARE_UF01.Q,
          dut.rw_reg.Q, dut.run_delay_reg.Q, dut.nextiv_ready_en_reg.Q, dut.hwrite_d1_reg.Q,
          dut.hready_resp_reg.Q, dut.deskey_unit.wr_ptr_reg_2.Q, dut.deskey_unit.wr_ptr_reg_1.Q,
          dut.deskey_unit.wr_ptr_reg_0.Q, dut.deskey_unit.ptr_reg_2.Q, dut.deskey_unit.ptr_reg_1.Q,
          dut.deskey_unit.ptr_reg_0.Q, dut.deskey_unit.fifo_mem_reg_5_31.Q, 
          dut.deskey_unit.fifo_mem_reg_5_30.Q, dut.deskey_unit.fifo_mem_reg_5_29.Q,
          dut.deskey_unit.fifo_mem_reg_5_28.Q, dut.deskey_unit.fifo_mem_reg_5_27.Q,
          dut.deskey_unit.fifo_mem_reg_5_26.Q, dut.deskey_unit.fifo_mem_reg_5_25.Q,
          dut.deskey_unit.fifo_mem_reg_5_23.Q, dut.deskey_unit.fifo_mem_reg_5_22.Q,
          dut.deskey_unit.fifo_mem_reg_5_21.Q, dut.deskey_unit.fifo_mem_reg_5_20.Q,
          dut.deskey_unit.fifo_mem_reg_5_19.Q, dut.deskey_unit.fifo_mem_reg_5_18.Q,
          dut.deskey_unit.fifo_mem_reg_5_17.Q, dut.deskey_unit.fifo_mem_reg_5_15.Q,
          dut.deskey_unit.fifo_mem_reg_5_14.Q, dut.deskey_unit.fifo_mem_reg_5_13.Q,
          dut.deskey_unit.fifo_mem_reg_5_12.Q, dut.deskey_unit.fifo_mem_reg_5_11.Q,
          dut.deskey_unit.fifo_mem_reg_5_10.Q, dut.deskey_unit.fifo_mem_reg_5_9.Q,
          dut.deskey_unit.fifo_mem_reg_5_7.Q, dut.deskey_unit.fifo_mem_reg_5_6.Q,
          dut.deskey_unit.fifo_mem_reg_5_5.Q, dut.deskey_unit.fifo_mem_reg_5_4.Q,
          dut.deskey_unit.fifo_mem_reg_5_3.Q, dut.deskey_unit.fifo_mem_reg_5_2.Q,
          dut.deskey_unit.fifo_mem_reg_5_1.Q, dut.deskey_unit.fifo_mem_reg_4_31.Q,
          dut.deskey_unit.fifo_mem_reg_4_30.Q, dut.deskey_unit.fifo_mem_reg_4_29.Q,
          dut.deskey_unit.fifo_mem_reg_4_28.Q, dut.deskey_unit.fifo_mem_reg_4_27.Q,
          dut.deskey_unit.fifo_mem_reg_4_26.Q, dut.deskey_unit.fifo_mem_reg_4_25.Q,
          dut.deskey_unit.fifo_mem_reg_4_23.Q, dut.deskey_unit.fifo_mem_reg_4_22.Q,
          dut.deskey_unit.fifo_mem_reg_4_21.Q, dut.deskey_unit.fifo_mem_reg_4_20.Q,
          dut.deskey_unit.fifo_mem_reg_4_19.Q, dut.deskey_unit.fifo_mem_reg_4_18.Q,
          dut.deskey_unit.fifo_mem_reg_4_17.Q, dut.deskey_unit.fifo_mem_reg_4_15.Q,
          dut.deskey_unit.fifo_mem_reg_4_14.Q, dut.deskey_unit.fifo_mem_reg_4_13.Q,
          dut.deskey_unit.fifo_mem_reg_4_12.Q, dut.deskey_unit.fifo_mem_reg_4_11.Q,
          dut.deskey_unit.fifo_mem_reg_4_10.Q, dut.deskey_unit.fifo_mem_reg_4_9.Q,
          dut.deskey_unit.fifo_mem_reg_4_7.Q, dut.deskey_unit.fifo_mem_reg_4_6.Q,
          dut.deskey_unit.fifo_mem_reg_4_5.Q, dut.deskey_unit.fifo_mem_reg_4_4.Q,
          dut.deskey_unit.fifo_mem_reg_4_3.Q, dut.deskey_unit.fifo_mem_reg_4_2.Q,
          dut.deskey_unit.fifo_mem_reg_4_1.Q, dut.deskey_unit.fifo_mem_reg_3_31.Q,
          dut.deskey_unit.fifo_mem_reg_3_30.Q, dut.deskey_unit.fifo_mem_reg_3_29.Q,
          dut.deskey_unit.fifo_mem_reg_3_28.Q, dut.deskey_unit.fifo_mem_reg_3_27.Q,
          dut.deskey_unit.fifo_mem_reg_3_26.Q, dut.deskey_unit.fifo_mem_reg_3_25.Q,
          dut.deskey_unit.fifo_mem_reg_3_23.Q, dut.deskey_unit.fifo_mem_reg_3_22.Q,
          dut.deskey_unit.fifo_mem_reg_3_21.Q, dut.deskey_unit.fifo_mem_reg_3_20.Q,
          dut.deskey_unit.fifo_mem_reg_3_19.Q, dut.deskey_unit.fifo_mem_reg_3_18.Q,
          dut.deskey_unit.fifo_mem_reg_3_17.Q, dut.deskey_unit.fifo_mem_reg_3_15.Q,
          dut.deskey_unit.fifo_mem_reg_3_14.Q, dut.deskey_unit.fifo_mem_reg_3_13.Q,
          dut.deskey_unit.fifo_mem_reg_3_12.Q, dut.deskey_unit.fifo_mem_reg_3_11.Q,
          dut.deskey_unit.fifo_mem_reg_3_10.Q, dut.deskey_unit.fifo_mem_reg_3_9.Q,
          dut.deskey_unit.fifo_mem_reg_3_7.Q, dut.deskey_unit.fifo_mem_reg_3_6.Q,
          dut.deskey_unit.fifo_mem_reg_3_5.Q, dut.deskey_unit.fifo_mem_reg_3_4.Q,
          dut.deskey_unit.fifo_mem_reg_3_3.Q, dut.deskey_unit.fifo_mem_reg_3_2.Q,
          dut.deskey_unit.fifo_mem_reg_3_1.Q, dut.deskey_unit.fifo_mem_reg_2_31.Q,
          dut.deskey_unit.fifo_mem_reg_2_30.Q, dut.deskey_unit.fifo_mem_reg_2_29.Q,
          dut.deskey_unit.fifo_mem_reg_2_28.Q, dut.deskey_unit.fifo_mem_reg_2_27.Q,
          dut.deskey_unit.fifo_mem_reg_2_26.Q, dut.deskey_unit.fifo_mem_reg_2_25.Q,
          dut.deskey_unit.fifo_mem_reg_2_23.Q, dut.deskey_unit.fifo_mem_reg_2_22.Q,
          dut.deskey_unit.fifo_mem_reg_2_21.Q, dut.deskey_unit.fifo_mem_reg_2_20.Q,
          dut.deskey_unit.fifo_mem_reg_2_19.Q, dut.deskey_unit.fifo_mem_reg_2_18.Q,
          dut.deskey_unit.fifo_mem_reg_2_17.Q, 1'b0 };

   event load_unload;
   always @ load_unload begin
      if (pattern != prev_pat) begin
         loads = 1;
         prev_pat = pattern;
         if ((verbose >= 2) && (pattern % report_interval == 0))
            $display("// %t : ...begin scan load for pattern %0d", $time, pattern);
         end
      else begin
         loads = loads + 1;
         if ((verbose >= 2) && (pattern % report_interval == 0))
            $display("// %t : ...begin scan load for pattern %0d, load %0d", $time, pattern, loads);
      end

      #0 PI[0] = 0; // hclk
      #0 PI[58] = 1'bX; // si0
      #0 PI[59] = 1'bX; // si1
      #0 PI[60] = 1'bX; // si2
      #0 PI[61] = 1'bX; // si3
      #0 PI[57] = 1; // Test_Se
      #0 PI[1] = 1; // POR
      #0 PI[56] = 1; // Test_Mode
      #0 PI[2] = 1; // hresetn
      #100;
      // end of load_unload preamble

      // gather current scan cell output bit values
      CHAINOUT[0] = (CHAINOUT0 ^ SHBEGM[0]) >> SHBEG;
      CHAINOUT[1] = (CHAINOUT1 ^ SHBEGM[1]) >> SHBEG;
      CHAINOUT[2] = (CHAINOUT2 ^ SHBEGM[2]) >> SHBEG;
      CHAINOUT[3] = (CHAINOUT3 ^ SHBEGM[3]) >> SHBEG;
      #0;

      // compare actual vs. expected values
      for (chain = 0; chain < 4; chain=chain + 1) begin
         UNL = UNLOAD[chain]; UNLM = UNLMSK[chain] & SERIALM; CHOUT = CHAINOUT[chain] ^ OUTINV[chain];
         if ((UNL&UNLM) !== (CHOUT&UNLM)) begin
            patp1 = pattern + lastpattern;  patm1 = patp1 - 1;
            if (lastpattern == 0) $display("\n// *** ERROR during scan pattern %0d (detected during load of pattern %0d), T=%t", patm1, patp1, $time );
            else                  $display("\n// *** ERROR during scan pattern %0d (detected during final pattern unload), T=%t", patm1, $time );
            for (bit = NSHIFTS+SHBEG; bit < LENMAX; bit=bit + 1) begin
               if ((UNL[bit]&UNLM[bit]) !== (CHOUT[bit]&UNLM[bit])) begin
                  $display("  %0d %0s %0d (exp=%b, got=%b)  // pin %0s, scan cell %0d",
                      patm1, CHAINnames[chain], bit, UNL[bit], CHOUT[bit], CHAINpins[chain], bit);
                  nofails = nofails + 1;
               end
            end
         end
      end
      #0;

      // force bits of scan chain 0
      LOADSH0 = (LOAD0 >> NSHIFTS) ^ INPINV[0];
      //force dut.desctrl_reg_4.TD = LOADSH0[0];
      force dut.desctrl_reg_3.TD = LOADSH0[1];
      force dut.desctrl_reg_2.TD = LOADSH0[2];
      force dut.desctrl_reg_1.TD = LOADSH0[3];
      force dut.desctrl_reg_0.TD = LOADSH0[4];
      force dut.des_cop_unit.flag_reg_1.TD = LOADSH0[5];
      force dut.des_cop_unit.flag_reg_0.TD = LOADSH0[6];
      force dut.des_cop_unit.din_valid_eins_reg.TD = LOADSH0[7];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_63.TD = LOADSH0[8];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_62.TD = LOADSH0[9];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_61.TD = LOADSH0[10];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_60.TD = LOADSH0[11];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_59.TD = LOADSH0[12];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_58.TD = LOADSH0[13];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_57.TD = LOADSH0[14];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_56.TD = LOADSH0[15];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_55.TD = LOADSH0[16];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_54.TD = LOADSH0[17];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_53.TD = LOADSH0[18];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_52.TD = LOADSH0[19];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_51.TD = LOADSH0[20];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_50.TD = LOADSH0[21];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_49.TD = LOADSH0[22];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_48.TD = LOADSH0[23];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_47.TD = LOADSH0[24];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_46.TD = LOADSH0[25];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_45.TD = LOADSH0[26];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_44.TD = LOADSH0[27];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_43.TD = LOADSH0[28];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_42.TD = LOADSH0[29];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_41.TD = LOADSH0[30];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_40.TD = LOADSH0[31];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_39.TD = LOADSH0[32];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_38.TD = LOADSH0[33];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_37.TD = LOADSH0[34];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_36.TD = LOADSH0[35];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_35.TD = LOADSH0[36];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_34.TD = LOADSH0[37];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_33.TD = LOADSH0[38];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_32.TD = LOADSH0[39];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_31.TD = LOADSH0[40];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_30.TD = LOADSH0[41];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_29.TD = LOADSH0[42];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_28.TD = LOADSH0[43];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_27.TD = LOADSH0[44];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_26.TD = LOADSH0[45];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_25.TD = LOADSH0[46];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_24.TD = LOADSH0[47];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_23.TD = LOADSH0[48];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_22.TD = LOADSH0[49];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_21.TD = LOADSH0[50];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_20.TD = LOADSH0[51];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_19.TD = LOADSH0[52];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_18.TD = LOADSH0[53];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_17.TD = LOADSH0[54];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_16.TD = LOADSH0[55];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_15.TD = LOADSH0[56];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_14.TD = LOADSH0[57];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_13.TD = LOADSH0[58];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_12.TD = LOADSH0[59];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_11.TD = LOADSH0[60];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_10.TD = LOADSH0[61];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_9.TD = LOADSH0[62];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_8.TD = LOADSH0[63];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_7.TD = LOADSH0[64];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_6.TD = LOADSH0[65];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_5.TD = LOADSH0[66];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_4.TD = LOADSH0[67];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_3.TD = LOADSH0[68];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_2.TD = LOADSH0[69];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_1.TD = LOADSH0[70];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_0.TD = LOADSH0[71];
      force dut.des_cop_unit.des_unit.u_tiny_des_round.clk_gate_obs.U1.TD = LOADSH0[72];
      force dut.des_cop_unit.des_unit.state_reg.TD = LOADSH0[73];
      force dut.des_cop_unit.des_unit.round_reg_3.TD = LOADSH0[74];
      force dut.des_cop_unit.des_unit.round_reg_2.TD = LOADSH0[75];
      force dut.des_cop_unit.des_unit.round_reg_1.TD = LOADSH0[76];
      force dut.des_cop_unit.des_unit.round_reg_0.TD = LOADSH0[77];
      force dut.des_cop_unit.des_unit.dout_valid_reg.TD = LOADSH0[78];
      force dut.data_in_reg_31.TD = LOADSH0[79];
      force dut.data_in_reg_30.TD = LOADSH0[80];
      force dut.data_in_reg_29.TD = LOADSH0[81];
      force dut.data_in_reg_28.TD = LOADSH0[82];
      force dut.data_in_reg_27.TD = LOADSH0[83];
      force dut.data_in_reg_26.TD = LOADSH0[84];
      force dut.data_in_reg_25.TD = LOADSH0[85];
      force dut.data_in_reg_24.TD = LOADSH0[86];
      force dut.data_in_reg_23.TD = LOADSH0[87];
      force dut.data_in_reg_22.TD = LOADSH0[88];
      force dut.data_in_reg_21.TD = LOADSH0[89];
      force dut.data_in_reg_20.TD = LOADSH0[90];
      force dut.data_in_reg_19.TD = LOADSH0[91];
      force dut.data_in_reg_18.TD = LOADSH0[92];
      force dut.data_in_reg_17.TD = LOADSH0[93];
      force dut.data_in_reg_16.TD = LOADSH0[94];
      force dut.data_in_reg_15.TD = LOADSH0[95];
      force dut.data_in_reg_14.TD = LOADSH0[96];
      force dut.data_in_reg_13.TD = LOADSH0[97];
      force dut.data_in_reg_12.TD = LOADSH0[98];
      force dut.data_in_reg_11.TD = LOADSH0[99];
      force dut.data_in_reg_10.TD = LOADSH0[100];
      force dut.data_in_reg_9.TD = LOADSH0[101];
      force dut.data_in_reg_8.TD = LOADSH0[102];
      force dut.data_in_reg_7.TD = LOADSH0[103];
      force dut.data_in_reg_6.TD = LOADSH0[104];
      force dut.data_in_reg_5.TD = LOADSH0[105];
      force dut.data_in_reg_4.TD = LOADSH0[106];
      force dut.data_in_reg_3.TD = LOADSH0[107];
      force dut.data_in_reg_2.TD = LOADSH0[108];
      force dut.data_in_reg_1.TD = LOADSH0[109];
      force dut.data_in_reg_0.TD = LOADSH0[110];
      force dut.clk_gate_obs.U1.TD = LOADSH0[111];

      // force bits of scan chain 1
      LOADSH1 = (LOAD1 >> NSHIFTS) ^ INPINV[1];
      //force dut.desiv_unit.fifo_mem_reg_0_28.TD = LOADSH1[1];
      force dut.desiv_unit.fifo_mem_reg_0_27.TD = LOADSH1[2];
      force dut.desiv_unit.fifo_mem_reg_0_26.TD = LOADSH1[3];
      force dut.desiv_unit.fifo_mem_reg_0_25.TD = LOADSH1[4];
      force dut.desiv_unit.fifo_mem_reg_0_24.TD = LOADSH1[5];
      force dut.desiv_unit.fifo_mem_reg_0_23.TD = LOADSH1[6];
      force dut.desiv_unit.fifo_mem_reg_0_22.TD = LOADSH1[7];
      force dut.desiv_unit.fifo_mem_reg_0_21.TD = LOADSH1[8];
      force dut.desiv_unit.fifo_mem_reg_0_20.TD = LOADSH1[9];
      force dut.desiv_unit.fifo_mem_reg_0_19.TD = LOADSH1[10];
      force dut.desiv_unit.fifo_mem_reg_0_18.TD = LOADSH1[11];
      force dut.desiv_unit.fifo_mem_reg_0_17.TD = LOADSH1[12];
      force dut.desiv_unit.fifo_mem_reg_0_16.TD = LOADSH1[13];
      force dut.desiv_unit.fifo_mem_reg_0_15.TD = LOADSH1[14];
      force dut.desiv_unit.fifo_mem_reg_0_14.TD = LOADSH1[15];
      force dut.desiv_unit.fifo_mem_reg_0_13.TD = LOADSH1[16];
      force dut.desiv_unit.fifo_mem_reg_0_12.TD = LOADSH1[17];
      force dut.desiv_unit.fifo_mem_reg_0_11.TD = LOADSH1[18];
      force dut.desiv_unit.fifo_mem_reg_0_10.TD = LOADSH1[19];
      force dut.desiv_unit.fifo_mem_reg_0_9.TD = LOADSH1[20];
      force dut.desiv_unit.fifo_mem_reg_0_8.TD = LOADSH1[21];
      force dut.desiv_unit.fifo_mem_reg_0_7.TD = LOADSH1[22];
      force dut.desiv_unit.fifo_mem_reg_0_6.TD = LOADSH1[23];
      force dut.desiv_unit.fifo_mem_reg_0_5.TD = LOADSH1[24];
      force dut.desiv_unit.fifo_mem_reg_0_4.TD = LOADSH1[25];
      force dut.desiv_unit.fifo_mem_reg_0_3.TD = LOADSH1[26];
      force dut.desiv_unit.fifo_mem_reg_0_2.TD = LOADSH1[27];
      force dut.desiv_unit.fifo_mem_reg_0_1.TD = LOADSH1[28];
      force dut.desiv_unit.fifo_mem_reg_0_0.TD = LOADSH1[29];
      force dut.desiv_unit.clk_gate_obs.U1.TD = LOADSH1[30];
      force dut.desiv_sel_reg.TD = LOADSH1[31];
      force dut.desiv_sel_d1_reg.TD = LOADSH1[32];
      force dut.desdat_unit.wr_ptr_reg.TD = LOADSH1[33];
      force dut.desdat_unit.rd_ptr_reg.TD = LOADSH1[34];
      force dut.desdat_unit.ptr_reg_1.TD = LOADSH1[35];
      force dut.desdat_unit.ptr_reg_0.TD = LOADSH1[36];
      force dut.desdat_unit.full_reg.TD = LOADSH1[37];
      force dut.desdat_unit.full_pulse_reg.TD = LOADSH1[38];
      force dut.desdat_unit.full_delay_reg.TD = LOADSH1[39];
      force dut.desdat_unit.fifo_mem_reg_1_31.TD = LOADSH1[40];
      force dut.desdat_unit.fifo_mem_reg_1_30.TD = LOADSH1[41];
      force dut.desdat_unit.fifo_mem_reg_1_29.TD = LOADSH1[42];
      force dut.desdat_unit.fifo_mem_reg_1_28.TD = LOADSH1[43];
      force dut.desdat_unit.fifo_mem_reg_1_27.TD = LOADSH1[44];
      force dut.desdat_unit.fifo_mem_reg_1_26.TD = LOADSH1[45];
      force dut.desdat_unit.fifo_mem_reg_1_25.TD = LOADSH1[46];
      force dut.desdat_unit.fifo_mem_reg_1_24.TD = LOADSH1[47];
      force dut.desdat_unit.fifo_mem_reg_1_23.TD = LOADSH1[48];
      force dut.desdat_unit.fifo_mem_reg_1_22.TD = LOADSH1[49];
      force dut.desdat_unit.fifo_mem_reg_1_21.TD = LOADSH1[50];
      force dut.desdat_unit.fifo_mem_reg_1_20.TD = LOADSH1[51];
      force dut.desdat_unit.fifo_mem_reg_1_19.TD = LOADSH1[52];
      force dut.desdat_unit.fifo_mem_reg_1_18.TD = LOADSH1[53];
      force dut.desdat_unit.fifo_mem_reg_1_17.TD = LOADSH1[54];
      force dut.desdat_unit.fifo_mem_reg_1_16.TD = LOADSH1[55];
      force dut.desdat_unit.fifo_mem_reg_1_15.TD = LOADSH1[56];
      force dut.desdat_unit.fifo_mem_reg_1_14.TD = LOADSH1[57];
      force dut.desdat_unit.fifo_mem_reg_1_13.TD = LOADSH1[58];
      force dut.desdat_unit.fifo_mem_reg_1_12.TD = LOADSH1[59];
      force dut.desdat_unit.fifo_mem_reg_1_11.TD = LOADSH1[60];
      force dut.desdat_unit.fifo_mem_reg_1_10.TD = LOADSH1[61];
      force dut.desdat_unit.fifo_mem_reg_1_9.TD = LOADSH1[62];
      force dut.desdat_unit.fifo_mem_reg_1_8.TD = LOADSH1[63];
      force dut.desdat_unit.fifo_mem_reg_1_7.TD = LOADSH1[64];
      force dut.desdat_unit.fifo_mem_reg_1_6.TD = LOADSH1[65];
      force dut.desdat_unit.fifo_mem_reg_1_5.TD = LOADSH1[66];
      force dut.desdat_unit.fifo_mem_reg_1_4.TD = LOADSH1[67];
      force dut.desdat_unit.fifo_mem_reg_1_3.TD = LOADSH1[68];
      force dut.desdat_unit.fifo_mem_reg_1_2.TD = LOADSH1[69];
      force dut.desdat_unit.fifo_mem_reg_1_1.TD = LOADSH1[70];
      force dut.desdat_unit.fifo_mem_reg_1_0.TD = LOADSH1[71];
      force dut.desdat_unit.fifo_mem_reg_0_31.TD = LOADSH1[72];
      force dut.desdat_unit.fifo_mem_reg_0_30.TD = LOADSH1[73];
      force dut.desdat_unit.fifo_mem_reg_0_29.TD = LOADSH1[74];
      force dut.desdat_unit.fifo_mem_reg_0_28.TD = LOADSH1[75];
      force dut.desdat_unit.fifo_mem_reg_0_27.TD = LOADSH1[76];
      force dut.desdat_unit.fifo_mem_reg_0_26.TD = LOADSH1[77];
      force dut.desdat_unit.fifo_mem_reg_0_25.TD = LOADSH1[78];
      force dut.desdat_unit.fifo_mem_reg_0_24.TD = LOADSH1[79];
      force dut.desdat_unit.fifo_mem_reg_0_23.TD = LOADSH1[80];
      force dut.desdat_unit.fifo_mem_reg_0_22.TD = LOADSH1[81];
      force dut.desdat_unit.fifo_mem_reg_0_21.TD = LOADSH1[82];
      force dut.desdat_unit.fifo_mem_reg_0_20.TD = LOADSH1[83];
      force dut.desdat_unit.fifo_mem_reg_0_19.TD = LOADSH1[84];
      force dut.desdat_unit.fifo_mem_reg_0_18.TD = LOADSH1[85];
      force dut.desdat_unit.fifo_mem_reg_0_17.TD = LOADSH1[86];
      force dut.desdat_unit.fifo_mem_reg_0_16.TD = LOADSH1[87];
      force dut.desdat_unit.fifo_mem_reg_0_15.TD = LOADSH1[88];
      force dut.desdat_unit.fifo_mem_reg_0_14.TD = LOADSH1[89];
      force dut.desdat_unit.fifo_mem_reg_0_13.TD = LOADSH1[90];
      force dut.desdat_unit.fifo_mem_reg_0_12.TD = LOADSH1[91];
      force dut.desdat_unit.fifo_mem_reg_0_11.TD = LOADSH1[92];
      force dut.desdat_unit.fifo_mem_reg_0_10.TD = LOADSH1[93];
      force dut.desdat_unit.fifo_mem_reg_0_9.TD = LOADSH1[94];
      force dut.desdat_unit.fifo_mem_reg_0_8.TD = LOADSH1[95];
      force dut.desdat_unit.fifo_mem_reg_0_7.TD = LOADSH1[96];
      force dut.desdat_unit.fifo_mem_reg_0_6.TD = LOADSH1[97];
      force dut.desdat_unit.fifo_mem_reg_0_5.TD = LOADSH1[98];
      force dut.desdat_unit.fifo_mem_reg_0_4.TD = LOADSH1[99];
      force dut.desdat_unit.fifo_mem_reg_0_3.TD = LOADSH1[100];
      force dut.desdat_unit.fifo_mem_reg_0_2.TD = LOADSH1[101];
      force dut.desdat_unit.fifo_mem_reg_0_1.TD = LOADSH1[102];
      force dut.desdat_unit.fifo_mem_reg_0_0.TD = LOADSH1[103];
      force dut.desdat_unit.clk_gate_obs.U1.TD = LOADSH1[104];
      force dut.desdat_sel_reg.TD = LOADSH1[105];
      force dut.desdat_sel_d1_reg.TD = LOADSH1[106];
      force dut.desctrl_sel_reg.TD = LOADSH1[107];
      force dut.desctrl_sel_d1_reg.TD = LOADSH1[108];
      force dut.desctrl_reg_7.TD = LOADSH1[109];
      force dut.desctrl_reg_6.TD = LOADSH1[110];
      force dut.desctrl_reg_5.TD = LOADSH1[111];

      // force bits of scan chain 2
      LOADSH2 = (LOAD2 >> NSHIFTS) ^ INPINV[2];
      //force dut.deskey_unit.fifo_mem_reg_2_15.TD = LOADSH2[1];
      force dut.deskey_unit.fifo_mem_reg_2_14.TD = LOADSH2[2];
      force dut.deskey_unit.fifo_mem_reg_2_13.TD = LOADSH2[3];
      force dut.deskey_unit.fifo_mem_reg_2_12.TD = LOADSH2[4];
      force dut.deskey_unit.fifo_mem_reg_2_11.TD = LOADSH2[5];
      force dut.deskey_unit.fifo_mem_reg_2_10.TD = LOADSH2[6];
      force dut.deskey_unit.fifo_mem_reg_2_9.TD = LOADSH2[7];
      force dut.deskey_unit.fifo_mem_reg_2_7.TD = LOADSH2[8];
      force dut.deskey_unit.fifo_mem_reg_2_6.TD = LOADSH2[9];
      force dut.deskey_unit.fifo_mem_reg_2_5.TD = LOADSH2[10];
      force dut.deskey_unit.fifo_mem_reg_2_4.TD = LOADSH2[11];
      force dut.deskey_unit.fifo_mem_reg_2_3.TD = LOADSH2[12];
      force dut.deskey_unit.fifo_mem_reg_2_2.TD = LOADSH2[13];
      force dut.deskey_unit.fifo_mem_reg_2_1.TD = LOADSH2[14];
      force dut.deskey_unit.fifo_mem_reg_1_31.TD = LOADSH2[15];
      force dut.deskey_unit.fifo_mem_reg_1_30.TD = LOADSH2[16];
      force dut.deskey_unit.fifo_mem_reg_1_29.TD = LOADSH2[17];
      force dut.deskey_unit.fifo_mem_reg_1_28.TD = LOADSH2[18];
      force dut.deskey_unit.fifo_mem_reg_1_27.TD = LOADSH2[19];
      force dut.deskey_unit.fifo_mem_reg_1_26.TD = LOADSH2[20];
      force dut.deskey_unit.fifo_mem_reg_1_25.TD = LOADSH2[21];
      force dut.deskey_unit.fifo_mem_reg_1_23.TD = LOADSH2[22];
      force dut.deskey_unit.fifo_mem_reg_1_22.TD = LOADSH2[23];
      force dut.deskey_unit.fifo_mem_reg_1_21.TD = LOADSH2[24];
      force dut.deskey_unit.fifo_mem_reg_1_20.TD = LOADSH2[25];
      force dut.deskey_unit.fifo_mem_reg_1_19.TD = LOADSH2[26];
      force dut.deskey_unit.fifo_mem_reg_1_18.TD = LOADSH2[27];
      force dut.deskey_unit.fifo_mem_reg_1_17.TD = LOADSH2[28];
      force dut.deskey_unit.fifo_mem_reg_1_15.TD = LOADSH2[29];
      force dut.deskey_unit.fifo_mem_reg_1_14.TD = LOADSH2[30];
      force dut.deskey_unit.fifo_mem_reg_1_13.TD = LOADSH2[31];
      force dut.deskey_unit.fifo_mem_reg_1_12.TD = LOADSH2[32];
      force dut.deskey_unit.fifo_mem_reg_1_11.TD = LOADSH2[33];
      force dut.deskey_unit.fifo_mem_reg_1_10.TD = LOADSH2[34];
      force dut.deskey_unit.fifo_mem_reg_1_9.TD = LOADSH2[35];
      force dut.deskey_unit.fifo_mem_reg_1_7.TD = LOADSH2[36];
      force dut.deskey_unit.fifo_mem_reg_1_6.TD = LOADSH2[37];
      force dut.deskey_unit.fifo_mem_reg_1_5.TD = LOADSH2[38];
      force dut.deskey_unit.fifo_mem_reg_1_4.TD = LOADSH2[39];
      force dut.deskey_unit.fifo_mem_reg_1_3.TD = LOADSH2[40];
      force dut.deskey_unit.fifo_mem_reg_1_2.TD = LOADSH2[41];
      force dut.deskey_unit.fifo_mem_reg_1_1.TD = LOADSH2[42];
      force dut.deskey_unit.fifo_mem_reg_0_31.TD = LOADSH2[43];
      force dut.deskey_unit.fifo_mem_reg_0_30.TD = LOADSH2[44];
      force dut.deskey_unit.fifo_mem_reg_0_29.TD = LOADSH2[45];
      force dut.deskey_unit.fifo_mem_reg_0_28.TD = LOADSH2[46];
      force dut.deskey_unit.fifo_mem_reg_0_27.TD = LOADSH2[47];
      force dut.deskey_unit.fifo_mem_reg_0_26.TD = LOADSH2[48];
      force dut.deskey_unit.fifo_mem_reg_0_25.TD = LOADSH2[49];
      force dut.deskey_unit.fifo_mem_reg_0_23.TD = LOADSH2[50];
      force dut.deskey_unit.fifo_mem_reg_0_22.TD = LOADSH2[51];
      force dut.deskey_unit.fifo_mem_reg_0_21.TD = LOADSH2[52];
      force dut.deskey_unit.fifo_mem_reg_0_20.TD = LOADSH2[53];
      force dut.deskey_unit.fifo_mem_reg_0_19.TD = LOADSH2[54];
      force dut.deskey_unit.fifo_mem_reg_0_18.TD = LOADSH2[55];
      force dut.deskey_unit.fifo_mem_reg_0_17.TD = LOADSH2[56];
      force dut.deskey_unit.fifo_mem_reg_0_15.TD = LOADSH2[57];
      force dut.deskey_unit.fifo_mem_reg_0_14.TD = LOADSH2[58];
      force dut.deskey_unit.fifo_mem_reg_0_13.TD = LOADSH2[59];
      force dut.deskey_unit.fifo_mem_reg_0_12.TD = LOADSH2[60];
      force dut.deskey_unit.fifo_mem_reg_0_11.TD = LOADSH2[61];
      force dut.deskey_unit.fifo_mem_reg_0_10.TD = LOADSH2[62];
      force dut.deskey_unit.fifo_mem_reg_0_9.TD = LOADSH2[63];
      force dut.deskey_unit.fifo_mem_reg_0_7.TD = LOADSH2[64];
      force dut.deskey_unit.fifo_mem_reg_0_6.TD = LOADSH2[65];
      force dut.deskey_unit.fifo_mem_reg_0_5.TD = LOADSH2[66];
      force dut.deskey_unit.fifo_mem_reg_0_4.TD = LOADSH2[67];
      force dut.deskey_unit.fifo_mem_reg_0_3.TD = LOADSH2[68];
      force dut.deskey_unit.fifo_mem_reg_0_2.TD = LOADSH2[69];
      force dut.deskey_unit.fifo_mem_reg_0_1.TD = LOADSH2[70];
      force dut.deskey_unit.clk_gate_obs.U1.TD = LOADSH2[71];
      force dut.deskey_sel_reg.TD = LOADSH2[72];
      force dut.deskey_sel_d1_reg.TD = LOADSH2[73];
      force dut.desiv_unit.wr_ptr_reg.TD = LOADSH2[74];
      force dut.desiv_unit.ptr_reg_1.TD = LOADSH2[75];
      force dut.desiv_unit.ptr_reg_0.TD = LOADSH2[76];
      force dut.desiv_unit.fifo_mem_reg_1_31.TD = LOADSH2[77];
      force dut.desiv_unit.fifo_mem_reg_1_30.TD = LOADSH2[78];
      force dut.desiv_unit.fifo_mem_reg_1_29.TD = LOADSH2[79];
      force dut.desiv_unit.fifo_mem_reg_1_28.TD = LOADSH2[80];
      force dut.desiv_unit.fifo_mem_reg_1_27.TD = LOADSH2[81];
      force dut.desiv_unit.fifo_mem_reg_1_26.TD = LOADSH2[82];
      force dut.desiv_unit.fifo_mem_reg_1_25.TD = LOADSH2[83];
      force dut.desiv_unit.fifo_mem_reg_1_24.TD = LOADSH2[84];
      force dut.desiv_unit.fifo_mem_reg_1_23.TD = LOADSH2[85];
      force dut.desiv_unit.fifo_mem_reg_1_22.TD = LOADSH2[86];
      force dut.desiv_unit.fifo_mem_reg_1_21.TD = LOADSH2[87];
      force dut.desiv_unit.fifo_mem_reg_1_20.TD = LOADSH2[88];
      force dut.desiv_unit.fifo_mem_reg_1_19.TD = LOADSH2[89];
      force dut.desiv_unit.fifo_mem_reg_1_18.TD = LOADSH2[90];
      force dut.desiv_unit.fifo_mem_reg_1_17.TD = LOADSH2[91];
      force dut.desiv_unit.fifo_mem_reg_1_16.TD = LOADSH2[92];
      force dut.desiv_unit.fifo_mem_reg_1_15.TD = LOADSH2[93];
      force dut.desiv_unit.fifo_mem_reg_1_14.TD = LOADSH2[94];
      force dut.desiv_unit.fifo_mem_reg_1_13.TD = LOADSH2[95];
      force dut.desiv_unit.fifo_mem_reg_1_12.TD = LOADSH2[96];
      force dut.desiv_unit.fifo_mem_reg_1_11.TD = LOADSH2[97];
      force dut.desiv_unit.fifo_mem_reg_1_10.TD = LOADSH2[98];
      force dut.desiv_unit.fifo_mem_reg_1_9.TD = LOADSH2[99];
      force dut.desiv_unit.fifo_mem_reg_1_8.TD = LOADSH2[100];
      force dut.desiv_unit.fifo_mem_reg_1_7.TD = LOADSH2[101];
      force dut.desiv_unit.fifo_mem_reg_1_6.TD = LOADSH2[102];
      force dut.desiv_unit.fifo_mem_reg_1_5.TD = LOADSH2[103];
      force dut.desiv_unit.fifo_mem_reg_1_4.TD = LOADSH2[104];
      force dut.desiv_unit.fifo_mem_reg_1_3.TD = LOADSH2[105];
      force dut.desiv_unit.fifo_mem_reg_1_2.TD = LOADSH2[106];
      force dut.desiv_unit.fifo_mem_reg_1_1.TD = LOADSH2[107];
      force dut.desiv_unit.fifo_mem_reg_1_0.TD = LOADSH2[108];
      force dut.desiv_unit.fifo_mem_reg_0_31.TD = LOADSH2[109];
      force dut.desiv_unit.fifo_mem_reg_0_30.TD = LOADSH2[110];
      force dut.desiv_unit.fifo_mem_reg_0_29.TD = LOADSH2[111];

      // force bits of scan chain 3
      LOADSH3 = (LOAD3 >> NSHIFTS) ^ INPINV[3];
      //force dut.u_des_spares_0.SPARE_UF03.TD = LOADSH3[1];
      force dut.u_des_spares_0.SPARE_UF01.TD = LOADSH3[2];
      force dut.rw_reg.TD = LOADSH3[3];
      force dut.run_delay_reg.TD = LOADSH3[4];
      force dut.nextiv_ready_en_reg.TD = LOADSH3[5];
      force dut.hwrite_d1_reg.TD = LOADSH3[6];
      force dut.hready_resp_reg.TD = LOADSH3[7];
      force dut.deskey_unit.wr_ptr_reg_2.TD = LOADSH3[8];
      force dut.deskey_unit.wr_ptr_reg_1.TD = LOADSH3[9];
      force dut.deskey_unit.wr_ptr_reg_0.TD = LOADSH3[10];
      force dut.deskey_unit.ptr_reg_2.TD = LOADSH3[11];
      force dut.deskey_unit.ptr_reg_1.TD = LOADSH3[12];
      force dut.deskey_unit.ptr_reg_0.TD = LOADSH3[13];
      force dut.deskey_unit.fifo_mem_reg_5_31.TD = LOADSH3[14];
      force dut.deskey_unit.fifo_mem_reg_5_30.TD = LOADSH3[15];
      force dut.deskey_unit.fifo_mem_reg_5_29.TD = LOADSH3[16];
      force dut.deskey_unit.fifo_mem_reg_5_28.TD = LOADSH3[17];
      force dut.deskey_unit.fifo_mem_reg_5_27.TD = LOADSH3[18];
      force dut.deskey_unit.fifo_mem_reg_5_26.TD = LOADSH3[19];
      force dut.deskey_unit.fifo_mem_reg_5_25.TD = LOADSH3[20];
      force dut.deskey_unit.fifo_mem_reg_5_23.TD = LOADSH3[21];
      force dut.deskey_unit.fifo_mem_reg_5_22.TD = LOADSH3[22];
      force dut.deskey_unit.fifo_mem_reg_5_21.TD = LOADSH3[23];
      force dut.deskey_unit.fifo_mem_reg_5_20.TD = LOADSH3[24];
      force dut.deskey_unit.fifo_mem_reg_5_19.TD = LOADSH3[25];
      force dut.deskey_unit.fifo_mem_reg_5_18.TD = LOADSH3[26];
      force dut.deskey_unit.fifo_mem_reg_5_17.TD = LOADSH3[27];
      force dut.deskey_unit.fifo_mem_reg_5_15.TD = LOADSH3[28];
      force dut.deskey_unit.fifo_mem_reg_5_14.TD = LOADSH3[29];
      force dut.deskey_unit.fifo_mem_reg_5_13.TD = LOADSH3[30];
      force dut.deskey_unit.fifo_mem_reg_5_12.TD = LOADSH3[31];
      force dut.deskey_unit.fifo_mem_reg_5_11.TD = LOADSH3[32];
      force dut.deskey_unit.fifo_mem_reg_5_10.TD = LOADSH3[33];
      force dut.deskey_unit.fifo_mem_reg_5_9.TD = LOADSH3[34];
      force dut.deskey_unit.fifo_mem_reg_5_7.TD = LOADSH3[35];
      force dut.deskey_unit.fifo_mem_reg_5_6.TD = LOADSH3[36];
      force dut.deskey_unit.fifo_mem_reg_5_5.TD = LOADSH3[37];
      force dut.deskey_unit.fifo_mem_reg_5_4.TD = LOADSH3[38];
      force dut.deskey_unit.fifo_mem_reg_5_3.TD = LOADSH3[39];
      force dut.deskey_unit.fifo_mem_reg_5_2.TD = LOADSH3[40];
      force dut.deskey_unit.fifo_mem_reg_5_1.TD = LOADSH3[41];
      force dut.deskey_unit.fifo_mem_reg_4_31.TD = LOADSH3[42];
      force dut.deskey_unit.fifo_mem_reg_4_30.TD = LOADSH3[43];
      force dut.deskey_unit.fifo_mem_reg_4_29.TD = LOADSH3[44];
      force dut.deskey_unit.fifo_mem_reg_4_28.TD = LOADSH3[45];
      force dut.deskey_unit.fifo_mem_reg_4_27.TD = LOADSH3[46];
      force dut.deskey_unit.fifo_mem_reg_4_26.TD = LOADSH3[47];
      force dut.deskey_unit.fifo_mem_reg_4_25.TD = LOADSH3[48];
      force dut.deskey_unit.fifo_mem_reg_4_23.TD = LOADSH3[49];
      force dut.deskey_unit.fifo_mem_reg_4_22.TD = LOADSH3[50];
      force dut.deskey_unit.fifo_mem_reg_4_21.TD = LOADSH3[51];
      force dut.deskey_unit.fifo_mem_reg_4_20.TD = LOADSH3[52];
      force dut.deskey_unit.fifo_mem_reg_4_19.TD = LOADSH3[53];
      force dut.deskey_unit.fifo_mem_reg_4_18.TD = LOADSH3[54];
      force dut.deskey_unit.fifo_mem_reg_4_17.TD = LOADSH3[55];
      force dut.deskey_unit.fifo_mem_reg_4_15.TD = LOADSH3[56];
      force dut.deskey_unit.fifo_mem_reg_4_14.TD = LOADSH3[57];
      force dut.deskey_unit.fifo_mem_reg_4_13.TD = LOADSH3[58];
      force dut.deskey_unit.fifo_mem_reg_4_12.TD = LOADSH3[59];
      force dut.deskey_unit.fifo_mem_reg_4_11.TD = LOADSH3[60];
      force dut.deskey_unit.fifo_mem_reg_4_10.TD = LOADSH3[61];
      force dut.deskey_unit.fifo_mem_reg_4_9.TD = LOADSH3[62];
      force dut.deskey_unit.fifo_mem_reg_4_7.TD = LOADSH3[63];
      force dut.deskey_unit.fifo_mem_reg_4_6.TD = LOADSH3[64];
      force dut.deskey_unit.fifo_mem_reg_4_5.TD = LOADSH3[65];
      force dut.deskey_unit.fifo_mem_reg_4_4.TD = LOADSH3[66];
      force dut.deskey_unit.fifo_mem_reg_4_3.TD = LOADSH3[67];
      force dut.deskey_unit.fifo_mem_reg_4_2.TD = LOADSH3[68];
      force dut.deskey_unit.fifo_mem_reg_4_1.TD = LOADSH3[69];
      force dut.deskey_unit.fifo_mem_reg_3_31.TD = LOADSH3[70];
      force dut.deskey_unit.fifo_mem_reg_3_30.TD = LOADSH3[71];
      force dut.deskey_unit.fifo_mem_reg_3_29.TD = LOADSH3[72];
      force dut.deskey_unit.fifo_mem_reg_3_28.TD = LOADSH3[73];
      force dut.deskey_unit.fifo_mem_reg_3_27.TD = LOADSH3[74];
      force dut.deskey_unit.fifo_mem_reg_3_26.TD = LOADSH3[75];
      force dut.deskey_unit.fifo_mem_reg_3_25.TD = LOADSH3[76];
      force dut.deskey_unit.fifo_mem_reg_3_23.TD = LOADSH3[77];
      force dut.deskey_unit.fifo_mem_reg_3_22.TD = LOADSH3[78];
      force dut.deskey_unit.fifo_mem_reg_3_21.TD = LOADSH3[79];
      force dut.deskey_unit.fifo_mem_reg_3_20.TD = LOADSH3[80];
      force dut.deskey_unit.fifo_mem_reg_3_19.TD = LOADSH3[81];
      force dut.deskey_unit.fifo_mem_reg_3_18.TD = LOADSH3[82];
      force dut.deskey_unit.fifo_mem_reg_3_17.TD = LOADSH3[83];
      force dut.deskey_unit.fifo_mem_reg_3_15.TD = LOADSH3[84];
      force dut.deskey_unit.fifo_mem_reg_3_14.TD = LOADSH3[85];
      force dut.deskey_unit.fifo_mem_reg_3_13.TD = LOADSH3[86];
      force dut.deskey_unit.fifo_mem_reg_3_12.TD = LOADSH3[87];
      force dut.deskey_unit.fifo_mem_reg_3_11.TD = LOADSH3[88];
      force dut.deskey_unit.fifo_mem_reg_3_10.TD = LOADSH3[89];
      force dut.deskey_unit.fifo_mem_reg_3_9.TD = LOADSH3[90];
      force dut.deskey_unit.fifo_mem_reg_3_7.TD = LOADSH3[91];
      force dut.deskey_unit.fifo_mem_reg_3_6.TD = LOADSH3[92];
      force dut.deskey_unit.fifo_mem_reg_3_5.TD = LOADSH3[93];
      force dut.deskey_unit.fifo_mem_reg_3_4.TD = LOADSH3[94];
      force dut.deskey_unit.fifo_mem_reg_3_3.TD = LOADSH3[95];
      force dut.deskey_unit.fifo_mem_reg_3_2.TD = LOADSH3[96];
      force dut.deskey_unit.fifo_mem_reg_3_1.TD = LOADSH3[97];
      force dut.deskey_unit.fifo_mem_reg_2_31.TD = LOADSH3[98];
      force dut.deskey_unit.fifo_mem_reg_2_30.TD = LOADSH3[99];
      force dut.deskey_unit.fifo_mem_reg_2_29.TD = LOADSH3[100];
      force dut.deskey_unit.fifo_mem_reg_2_28.TD = LOADSH3[101];
      force dut.deskey_unit.fifo_mem_reg_2_27.TD = LOADSH3[102];
      force dut.deskey_unit.fifo_mem_reg_2_26.TD = LOADSH3[103];
      force dut.deskey_unit.fifo_mem_reg_2_25.TD = LOADSH3[104];
      force dut.deskey_unit.fifo_mem_reg_2_23.TD = LOADSH3[105];
      force dut.deskey_unit.fifo_mem_reg_2_22.TD = LOADSH3[106];
      force dut.deskey_unit.fifo_mem_reg_2_21.TD = LOADSH3[107];
      force dut.deskey_unit.fifo_mem_reg_2_20.TD = LOADSH3[108];
      force dut.deskey_unit.fifo_mem_reg_2_19.TD = LOADSH3[109];
      force dut.deskey_unit.fifo_mem_reg_2_18.TD = LOADSH3[110];
      force dut.deskey_unit.fifo_mem_reg_2_17.TD = LOADSH3[111];
      #0;

      // apply single shift pulse with force's in place
      bit = LENMAX - NSHIFTS - 1;
      shift;

      // release bits of scan chain 0
      //release dut.desctrl_reg_4.TD;
      release dut.desctrl_reg_3.TD;
      release dut.desctrl_reg_2.TD;
      release dut.desctrl_reg_1.TD;
      release dut.desctrl_reg_0.TD;
      release dut.des_cop_unit.flag_reg_1.TD;
      release dut.des_cop_unit.flag_reg_0.TD;
      release dut.des_cop_unit.din_valid_eins_reg.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_63.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_62.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_61.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_60.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_59.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_58.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_57.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_56.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_55.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_54.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_53.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_52.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_51.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_50.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_49.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_48.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_47.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_46.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_45.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_44.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_43.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_42.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_41.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_40.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_39.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_38.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_37.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_36.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_35.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_34.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_33.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_32.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_31.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_30.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_29.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_28.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_27.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_26.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_25.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_24.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_23.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_22.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_21.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_20.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_19.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_18.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_17.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_16.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_15.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_14.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_13.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_12.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_11.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_10.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_9.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_8.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_7.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_6.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_5.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_4.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_3.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_2.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_1.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.dout_reg_0.TD;
      release dut.des_cop_unit.des_unit.u_tiny_des_round.clk_gate_obs.U1.TD;
      release dut.des_cop_unit.des_unit.state_reg.TD;
      release dut.des_cop_unit.des_unit.round_reg_3.TD;
      release dut.des_cop_unit.des_unit.round_reg_2.TD;
      release dut.des_cop_unit.des_unit.round_reg_1.TD;
      release dut.des_cop_unit.des_unit.round_reg_0.TD;
      release dut.des_cop_unit.des_unit.dout_valid_reg.TD;
      release dut.data_in_reg_31.TD;
      release dut.data_in_reg_30.TD;
      release dut.data_in_reg_29.TD;
      release dut.data_in_reg_28.TD;
      release dut.data_in_reg_27.TD;
      release dut.data_in_reg_26.TD;
      release dut.data_in_reg_25.TD;
      release dut.data_in_reg_24.TD;
      release dut.data_in_reg_23.TD;
      release dut.data_in_reg_22.TD;
      release dut.data_in_reg_21.TD;
      release dut.data_in_reg_20.TD;
      release dut.data_in_reg_19.TD;
      release dut.data_in_reg_18.TD;
      release dut.data_in_reg_17.TD;
      release dut.data_in_reg_16.TD;
      release dut.data_in_reg_15.TD;
      release dut.data_in_reg_14.TD;
      release dut.data_in_reg_13.TD;
      release dut.data_in_reg_12.TD;
      release dut.data_in_reg_11.TD;
      release dut.data_in_reg_10.TD;
      release dut.data_in_reg_9.TD;
      release dut.data_in_reg_8.TD;
      release dut.data_in_reg_7.TD;
      release dut.data_in_reg_6.TD;
      release dut.data_in_reg_5.TD;
      release dut.data_in_reg_4.TD;
      release dut.data_in_reg_3.TD;
      release dut.data_in_reg_2.TD;
      release dut.data_in_reg_1.TD;
      release dut.data_in_reg_0.TD;
      release dut.clk_gate_obs.U1.TD;

      // release bits of scan chain 1
      //release dut.desiv_unit.fifo_mem_reg_0_28.TD;
      release dut.desiv_unit.fifo_mem_reg_0_27.TD;
      release dut.desiv_unit.fifo_mem_reg_0_26.TD;
      release dut.desiv_unit.fifo_mem_reg_0_25.TD;
      release dut.desiv_unit.fifo_mem_reg_0_24.TD;
      release dut.desiv_unit.fifo_mem_reg_0_23.TD;
      release dut.desiv_unit.fifo_mem_reg_0_22.TD;
      release dut.desiv_unit.fifo_mem_reg_0_21.TD;
      release dut.desiv_unit.fifo_mem_reg_0_20.TD;
      release dut.desiv_unit.fifo_mem_reg_0_19.TD;
      release dut.desiv_unit.fifo_mem_reg_0_18.TD;
      release dut.desiv_unit.fifo_mem_reg_0_17.TD;
      release dut.desiv_unit.fifo_mem_reg_0_16.TD;
      release dut.desiv_unit.fifo_mem_reg_0_15.TD;
      release dut.desiv_unit.fifo_mem_reg_0_14.TD;
      release dut.desiv_unit.fifo_mem_reg_0_13.TD;
      release dut.desiv_unit.fifo_mem_reg_0_12.TD;
      release dut.desiv_unit.fifo_mem_reg_0_11.TD;
      release dut.desiv_unit.fifo_mem_reg_0_10.TD;
      release dut.desiv_unit.fifo_mem_reg_0_9.TD;
      release dut.desiv_unit.fifo_mem_reg_0_8.TD;
      release dut.desiv_unit.fifo_mem_reg_0_7.TD;
      release dut.desiv_unit.fifo_mem_reg_0_6.TD;
      release dut.desiv_unit.fifo_mem_reg_0_5.TD;
      release dut.desiv_unit.fifo_mem_reg_0_4.TD;
      release dut.desiv_unit.fifo_mem_reg_0_3.TD;
      release dut.desiv_unit.fifo_mem_reg_0_2.TD;
      release dut.desiv_unit.fifo_mem_reg_0_1.TD;
      release dut.desiv_unit.fifo_mem_reg_0_0.TD;
      release dut.desiv_unit.clk_gate_obs.U1.TD;
      release dut.desiv_sel_reg.TD;
      release dut.desiv_sel_d1_reg.TD;
      release dut.desdat_unit.wr_ptr_reg.TD;
      release dut.desdat_unit.rd_ptr_reg.TD;
      release dut.desdat_unit.ptr_reg_1.TD;
      release dut.desdat_unit.ptr_reg_0.TD;
      release dut.desdat_unit.full_reg.TD;
      release dut.desdat_unit.full_pulse_reg.TD;
      release dut.desdat_unit.full_delay_reg.TD;
      release dut.desdat_unit.fifo_mem_reg_1_31.TD;
      release dut.desdat_unit.fifo_mem_reg_1_30.TD;
      release dut.desdat_unit.fifo_mem_reg_1_29.TD;
      release dut.desdat_unit.fifo_mem_reg_1_28.TD;
      release dut.desdat_unit.fifo_mem_reg_1_27.TD;
      release dut.desdat_unit.fifo_mem_reg_1_26.TD;
      release dut.desdat_unit.fifo_mem_reg_1_25.TD;
      release dut.desdat_unit.fifo_mem_reg_1_24.TD;
      release dut.desdat_unit.fifo_mem_reg_1_23.TD;
      release dut.desdat_unit.fifo_mem_reg_1_22.TD;
      release dut.desdat_unit.fifo_mem_reg_1_21.TD;
      release dut.desdat_unit.fifo_mem_reg_1_20.TD;
      release dut.desdat_unit.fifo_mem_reg_1_19.TD;
      release dut.desdat_unit.fifo_mem_reg_1_18.TD;
      release dut.desdat_unit.fifo_mem_reg_1_17.TD;
      release dut.desdat_unit.fifo_mem_reg_1_16.TD;
      release dut.desdat_unit.fifo_mem_reg_1_15.TD;
      release dut.desdat_unit.fifo_mem_reg_1_14.TD;
      release dut.desdat_unit.fifo_mem_reg_1_13.TD;
      release dut.desdat_unit.fifo_mem_reg_1_12.TD;
      release dut.desdat_unit.fifo_mem_reg_1_11.TD;
      release dut.desdat_unit.fifo_mem_reg_1_10.TD;
      release dut.desdat_unit.fifo_mem_reg_1_9.TD;
      release dut.desdat_unit.fifo_mem_reg_1_8.TD;
      release dut.desdat_unit.fifo_mem_reg_1_7.TD;
      release dut.desdat_unit.fifo_mem_reg_1_6.TD;
      release dut.desdat_unit.fifo_mem_reg_1_5.TD;
      release dut.desdat_unit.fifo_mem_reg_1_4.TD;
      release dut.desdat_unit.fifo_mem_reg_1_3.TD;
      release dut.desdat_unit.fifo_mem_reg_1_2.TD;
      release dut.desdat_unit.fifo_mem_reg_1_1.TD;
      release dut.desdat_unit.fifo_mem_reg_1_0.TD;
      release dut.desdat_unit.fifo_mem_reg_0_31.TD;
      release dut.desdat_unit.fifo_mem_reg_0_30.TD;
      release dut.desdat_unit.fifo_mem_reg_0_29.TD;
      release dut.desdat_unit.fifo_mem_reg_0_28.TD;
      release dut.desdat_unit.fifo_mem_reg_0_27.TD;
      release dut.desdat_unit.fifo_mem_reg_0_26.TD;
      release dut.desdat_unit.fifo_mem_reg_0_25.TD;
      release dut.desdat_unit.fifo_mem_reg_0_24.TD;
      release dut.desdat_unit.fifo_mem_reg_0_23.TD;
      release dut.desdat_unit.fifo_mem_reg_0_22.TD;
      release dut.desdat_unit.fifo_mem_reg_0_21.TD;
      release dut.desdat_unit.fifo_mem_reg_0_20.TD;
      release dut.desdat_unit.fifo_mem_reg_0_19.TD;
      release dut.desdat_unit.fifo_mem_reg_0_18.TD;
      release dut.desdat_unit.fifo_mem_reg_0_17.TD;
      release dut.desdat_unit.fifo_mem_reg_0_16.TD;
      release dut.desdat_unit.fifo_mem_reg_0_15.TD;
      release dut.desdat_unit.fifo_mem_reg_0_14.TD;
      release dut.desdat_unit.fifo_mem_reg_0_13.TD;
      release dut.desdat_unit.fifo_mem_reg_0_12.TD;
      release dut.desdat_unit.fifo_mem_reg_0_11.TD;
      release dut.desdat_unit.fifo_mem_reg_0_10.TD;
      release dut.desdat_unit.fifo_mem_reg_0_9.TD;
      release dut.desdat_unit.fifo_mem_reg_0_8.TD;
      release dut.desdat_unit.fifo_mem_reg_0_7.TD;
      release dut.desdat_unit.fifo_mem_reg_0_6.TD;
      release dut.desdat_unit.fifo_mem_reg_0_5.TD;
      release dut.desdat_unit.fifo_mem_reg_0_4.TD;
      release dut.desdat_unit.fifo_mem_reg_0_3.TD;
      release dut.desdat_unit.fifo_mem_reg_0_2.TD;
      release dut.desdat_unit.fifo_mem_reg_0_1.TD;
      release dut.desdat_unit.fifo_mem_reg_0_0.TD;
      release dut.desdat_unit.clk_gate_obs.U1.TD;
      release dut.desdat_sel_reg.TD;
      release dut.desdat_sel_d1_reg.TD;
      release dut.desctrl_sel_reg.TD;
      release dut.desctrl_sel_d1_reg.TD;
      release dut.desctrl_reg_7.TD;
      release dut.desctrl_reg_6.TD;
      release dut.desctrl_reg_5.TD;

      // release bits of scan chain 2
      //release dut.deskey_unit.fifo_mem_reg_2_15.TD;
      release dut.deskey_unit.fifo_mem_reg_2_14.TD;
      release dut.deskey_unit.fifo_mem_reg_2_13.TD;
      release dut.deskey_unit.fifo_mem_reg_2_12.TD;
      release dut.deskey_unit.fifo_mem_reg_2_11.TD;
      release dut.deskey_unit.fifo_mem_reg_2_10.TD;
      release dut.deskey_unit.fifo_mem_reg_2_9.TD;
      release dut.deskey_unit.fifo_mem_reg_2_7.TD;
      release dut.deskey_unit.fifo_mem_reg_2_6.TD;
      release dut.deskey_unit.fifo_mem_reg_2_5.TD;
      release dut.deskey_unit.fifo_mem_reg_2_4.TD;
      release dut.deskey_unit.fifo_mem_reg_2_3.TD;
      release dut.deskey_unit.fifo_mem_reg_2_2.TD;
      release dut.deskey_unit.fifo_mem_reg_2_1.TD;
      release dut.deskey_unit.fifo_mem_reg_1_31.TD;
      release dut.deskey_unit.fifo_mem_reg_1_30.TD;
      release dut.deskey_unit.fifo_mem_reg_1_29.TD;
      release dut.deskey_unit.fifo_mem_reg_1_28.TD;
      release dut.deskey_unit.fifo_mem_reg_1_27.TD;
      release dut.deskey_unit.fifo_mem_reg_1_26.TD;
      release dut.deskey_unit.fifo_mem_reg_1_25.TD;
      release dut.deskey_unit.fifo_mem_reg_1_23.TD;
      release dut.deskey_unit.fifo_mem_reg_1_22.TD;
      release dut.deskey_unit.fifo_mem_reg_1_21.TD;
      release dut.deskey_unit.fifo_mem_reg_1_20.TD;
      release dut.deskey_unit.fifo_mem_reg_1_19.TD;
      release dut.deskey_unit.fifo_mem_reg_1_18.TD;
      release dut.deskey_unit.fifo_mem_reg_1_17.TD;
      release dut.deskey_unit.fifo_mem_reg_1_15.TD;
      release dut.deskey_unit.fifo_mem_reg_1_14.TD;
      release dut.deskey_unit.fifo_mem_reg_1_13.TD;
      release dut.deskey_unit.fifo_mem_reg_1_12.TD;
      release dut.deskey_unit.fifo_mem_reg_1_11.TD;
      release dut.deskey_unit.fifo_mem_reg_1_10.TD;
      release dut.deskey_unit.fifo_mem_reg_1_9.TD;
      release dut.deskey_unit.fifo_mem_reg_1_7.TD;
      release dut.deskey_unit.fifo_mem_reg_1_6.TD;
      release dut.deskey_unit.fifo_mem_reg_1_5.TD;
      release dut.deskey_unit.fifo_mem_reg_1_4.TD;
      release dut.deskey_unit.fifo_mem_reg_1_3.TD;
      release dut.deskey_unit.fifo_mem_reg_1_2.TD;
      release dut.deskey_unit.fifo_mem_reg_1_1.TD;
      release dut.deskey_unit.fifo_mem_reg_0_31.TD;
      release dut.deskey_unit.fifo_mem_reg_0_30.TD;
      release dut.deskey_unit.fifo_mem_reg_0_29.TD;
      release dut.deskey_unit.fifo_mem_reg_0_28.TD;
      release dut.deskey_unit.fifo_mem_reg_0_27.TD;
      release dut.deskey_unit.fifo_mem_reg_0_26.TD;
      release dut.deskey_unit.fifo_mem_reg_0_25.TD;
      release dut.deskey_unit.fifo_mem_reg_0_23.TD;
      release dut.deskey_unit.fifo_mem_reg_0_22.TD;
      release dut.deskey_unit.fifo_mem_reg_0_21.TD;
      release dut.deskey_unit.fifo_mem_reg_0_20.TD;
      release dut.deskey_unit.fifo_mem_reg_0_19.TD;
      release dut.deskey_unit.fifo_mem_reg_0_18.TD;
      release dut.deskey_unit.fifo_mem_reg_0_17.TD;
      release dut.deskey_unit.fifo_mem_reg_0_15.TD;
      release dut.deskey_unit.fifo_mem_reg_0_14.TD;
      release dut.deskey_unit.fifo_mem_reg_0_13.TD;
      release dut.deskey_unit.fifo_mem_reg_0_12.TD;
      release dut.deskey_unit.fifo_mem_reg_0_11.TD;
      release dut.deskey_unit.fifo_mem_reg_0_10.TD;
      release dut.deskey_unit.fifo_mem_reg_0_9.TD;
      release dut.deskey_unit.fifo_mem_reg_0_7.TD;
      release dut.deskey_unit.fifo_mem_reg_0_6.TD;
      release dut.deskey_unit.fifo_mem_reg_0_5.TD;
      release dut.deskey_unit.fifo_mem_reg_0_4.TD;
      release dut.deskey_unit.fifo_mem_reg_0_3.TD;
      release dut.deskey_unit.fifo_mem_reg_0_2.TD;
      release dut.deskey_unit.fifo_mem_reg_0_1.TD;
      release dut.deskey_unit.clk_gate_obs.U1.TD;
      release dut.deskey_sel_reg.TD;
      release dut.deskey_sel_d1_reg.TD;
      release dut.desiv_unit.wr_ptr_reg.TD;
      release dut.desiv_unit.ptr_reg_1.TD;
      release dut.desiv_unit.ptr_reg_0.TD;
      release dut.desiv_unit.fifo_mem_reg_1_31.TD;
      release dut.desiv_unit.fifo_mem_reg_1_30.TD;
      release dut.desiv_unit.fifo_mem_reg_1_29.TD;
      release dut.desiv_unit.fifo_mem_reg_1_28.TD;
      release dut.desiv_unit.fifo_mem_reg_1_27.TD;
      release dut.desiv_unit.fifo_mem_reg_1_26.TD;
      release dut.desiv_unit.fifo_mem_reg_1_25.TD;
      release dut.desiv_unit.fifo_mem_reg_1_24.TD;
      release dut.desiv_unit.fifo_mem_reg_1_23.TD;
      release dut.desiv_unit.fifo_mem_reg_1_22.TD;
      release dut.desiv_unit.fifo_mem_reg_1_21.TD;
      release dut.desiv_unit.fifo_mem_reg_1_20.TD;
      release dut.desiv_unit.fifo_mem_reg_1_19.TD;
      release dut.desiv_unit.fifo_mem_reg_1_18.TD;
      release dut.desiv_unit.fifo_mem_reg_1_17.TD;
      release dut.desiv_unit.fifo_mem_reg_1_16.TD;
      release dut.desiv_unit.fifo_mem_reg_1_15.TD;
      release dut.desiv_unit.fifo_mem_reg_1_14.TD;
      release dut.desiv_unit.fifo_mem_reg_1_13.TD;
      release dut.desiv_unit.fifo_mem_reg_1_12.TD;
      release dut.desiv_unit.fifo_mem_reg_1_11.TD;
      release dut.desiv_unit.fifo_mem_reg_1_10.TD;
      release dut.desiv_unit.fifo_mem_reg_1_9.TD;
      release dut.desiv_unit.fifo_mem_reg_1_8.TD;
      release dut.desiv_unit.fifo_mem_reg_1_7.TD;
      release dut.desiv_unit.fifo_mem_reg_1_6.TD;
      release dut.desiv_unit.fifo_mem_reg_1_5.TD;
      release dut.desiv_unit.fifo_mem_reg_1_4.TD;
      release dut.desiv_unit.fifo_mem_reg_1_3.TD;
      release dut.desiv_unit.fifo_mem_reg_1_2.TD;
      release dut.desiv_unit.fifo_mem_reg_1_1.TD;
      release dut.desiv_unit.fifo_mem_reg_1_0.TD;
      release dut.desiv_unit.fifo_mem_reg_0_31.TD;
      release dut.desiv_unit.fifo_mem_reg_0_30.TD;
      release dut.desiv_unit.fifo_mem_reg_0_29.TD;

      // release bits of scan chain 3
      //release dut.u_des_spares_0.SPARE_UF03.TD;
      release dut.u_des_spares_0.SPARE_UF01.TD;
      release dut.rw_reg.TD;
      release dut.run_delay_reg.TD;
      release dut.nextiv_ready_en_reg.TD;
      release dut.hwrite_d1_reg.TD;
      release dut.hready_resp_reg.TD;
      release dut.deskey_unit.wr_ptr_reg_2.TD;
      release dut.deskey_unit.wr_ptr_reg_1.TD;
      release dut.deskey_unit.wr_ptr_reg_0.TD;
      release dut.deskey_unit.ptr_reg_2.TD;
      release dut.deskey_unit.ptr_reg_1.TD;
      release dut.deskey_unit.ptr_reg_0.TD;
      release dut.deskey_unit.fifo_mem_reg_5_31.TD;
      release dut.deskey_unit.fifo_mem_reg_5_30.TD;
      release dut.deskey_unit.fifo_mem_reg_5_29.TD;
      release dut.deskey_unit.fifo_mem_reg_5_28.TD;
      release dut.deskey_unit.fifo_mem_reg_5_27.TD;
      release dut.deskey_unit.fifo_mem_reg_5_26.TD;
      release dut.deskey_unit.fifo_mem_reg_5_25.TD;
      release dut.deskey_unit.fifo_mem_reg_5_23.TD;
      release dut.deskey_unit.fifo_mem_reg_5_22.TD;
      release dut.deskey_unit.fifo_mem_reg_5_21.TD;
      release dut.deskey_unit.fifo_mem_reg_5_20.TD;
      release dut.deskey_unit.fifo_mem_reg_5_19.TD;
      release dut.deskey_unit.fifo_mem_reg_5_18.TD;
      release dut.deskey_unit.fifo_mem_reg_5_17.TD;
      release dut.deskey_unit.fifo_mem_reg_5_15.TD;
      release dut.deskey_unit.fifo_mem_reg_5_14.TD;
      release dut.deskey_unit.fifo_mem_reg_5_13.TD;
      release dut.deskey_unit.fifo_mem_reg_5_12.TD;
      release dut.deskey_unit.fifo_mem_reg_5_11.TD;
      release dut.deskey_unit.fifo_mem_reg_5_10.TD;
      release dut.deskey_unit.fifo_mem_reg_5_9.TD;
      release dut.deskey_unit.fifo_mem_reg_5_7.TD;
      release dut.deskey_unit.fifo_mem_reg_5_6.TD;
      release dut.deskey_unit.fifo_mem_reg_5_5.TD;
      release dut.deskey_unit.fifo_mem_reg_5_4.TD;
      release dut.deskey_unit.fifo_mem_reg_5_3.TD;
      release dut.deskey_unit.fifo_mem_reg_5_2.TD;
      release dut.deskey_unit.fifo_mem_reg_5_1.TD;
      release dut.deskey_unit.fifo_mem_reg_4_31.TD;
      release dut.deskey_unit.fifo_mem_reg_4_30.TD;
      release dut.deskey_unit.fifo_mem_reg_4_29.TD;
      release dut.deskey_unit.fifo_mem_reg_4_28.TD;
      release dut.deskey_unit.fifo_mem_reg_4_27.TD;
      release dut.deskey_unit.fifo_mem_reg_4_26.TD;
      release dut.deskey_unit.fifo_mem_reg_4_25.TD;
      release dut.deskey_unit.fifo_mem_reg_4_23.TD;
      release dut.deskey_unit.fifo_mem_reg_4_22.TD;
      release dut.deskey_unit.fifo_mem_reg_4_21.TD;
      release dut.deskey_unit.fifo_mem_reg_4_20.TD;
      release dut.deskey_unit.fifo_mem_reg_4_19.TD;
      release dut.deskey_unit.fifo_mem_reg_4_18.TD;
      release dut.deskey_unit.fifo_mem_reg_4_17.TD;
      release dut.deskey_unit.fifo_mem_reg_4_15.TD;
      release dut.deskey_unit.fifo_mem_reg_4_14.TD;
      release dut.deskey_unit.fifo_mem_reg_4_13.TD;
      release dut.deskey_unit.fifo_mem_reg_4_12.TD;
      release dut.deskey_unit.fifo_mem_reg_4_11.TD;
      release dut.deskey_unit.fifo_mem_reg_4_10.TD;
      release dut.deskey_unit.fifo_mem_reg_4_9.TD;
      release dut.deskey_unit.fifo_mem_reg_4_7.TD;
      release dut.deskey_unit.fifo_mem_reg_4_6.TD;
      release dut.deskey_unit.fifo_mem_reg_4_5.TD;
      release dut.deskey_unit.fifo_mem_reg_4_4.TD;
      release dut.deskey_unit.fifo_mem_reg_4_3.TD;
      release dut.deskey_unit.fifo_mem_reg_4_2.TD;
      release dut.deskey_unit.fifo_mem_reg_4_1.TD;
      release dut.deskey_unit.fifo_mem_reg_3_31.TD;
      release dut.deskey_unit.fifo_mem_reg_3_30.TD;
      release dut.deskey_unit.fifo_mem_reg_3_29.TD;
      release dut.deskey_unit.fifo_mem_reg_3_28.TD;
      release dut.deskey_unit.fifo_mem_reg_3_27.TD;
      release dut.deskey_unit.fifo_mem_reg_3_26.TD;
      release dut.deskey_unit.fifo_mem_reg_3_25.TD;
      release dut.deskey_unit.fifo_mem_reg_3_23.TD;
      release dut.deskey_unit.fifo_mem_reg_3_22.TD;
      release dut.deskey_unit.fifo_mem_reg_3_21.TD;
      release dut.deskey_unit.fifo_mem_reg_3_20.TD;
      release dut.deskey_unit.fifo_mem_reg_3_19.TD;
      release dut.deskey_unit.fifo_mem_reg_3_18.TD;
      release dut.deskey_unit.fifo_mem_reg_3_17.TD;
      release dut.deskey_unit.fifo_mem_reg_3_15.TD;
      release dut.deskey_unit.fifo_mem_reg_3_14.TD;
      release dut.deskey_unit.fifo_mem_reg_3_13.TD;
      release dut.deskey_unit.fifo_mem_reg_3_12.TD;
      release dut.deskey_unit.fifo_mem_reg_3_11.TD;
      release dut.deskey_unit.fifo_mem_reg_3_10.TD;
      release dut.deskey_unit.fifo_mem_reg_3_9.TD;
      release dut.deskey_unit.fifo_mem_reg_3_7.TD;
      release dut.deskey_unit.fifo_mem_reg_3_6.TD;
      release dut.deskey_unit.fifo_mem_reg_3_5.TD;
      release dut.deskey_unit.fifo_mem_reg_3_4.TD;
      release dut.deskey_unit.fifo_mem_reg_3_3.TD;
      release dut.deskey_unit.fifo_mem_reg_3_2.TD;
      release dut.deskey_unit.fifo_mem_reg_3_1.TD;
      release dut.deskey_unit.fifo_mem_reg_2_31.TD;
      release dut.deskey_unit.fifo_mem_reg_2_30.TD;
      release dut.deskey_unit.fifo_mem_reg_2_29.TD;
      release dut.deskey_unit.fifo_mem_reg_2_28.TD;
      release dut.deskey_unit.fifo_mem_reg_2_27.TD;
      release dut.deskey_unit.fifo_mem_reg_2_26.TD;
      release dut.deskey_unit.fifo_mem_reg_2_25.TD;
      release dut.deskey_unit.fifo_mem_reg_2_23.TD;
      release dut.deskey_unit.fifo_mem_reg_2_22.TD;
      release dut.deskey_unit.fifo_mem_reg_2_21.TD;
      release dut.deskey_unit.fifo_mem_reg_2_20.TD;
      release dut.deskey_unit.fifo_mem_reg_2_19.TD;
      release dut.deskey_unit.fifo_mem_reg_2_18.TD;
      release dut.deskey_unit.fifo_mem_reg_2_17.TD;
      #0;

      // handle potential of last N bits shifted serially
      if (NSHIFTS > SHEND) begin
         bit = LENMAX-NSHIFTS; multiple_shift;
      end
   end

   `ifdef tmax_serial_timing
      parameter load_delay = 11300; // equivalent serial simulation load_unload time advance
   `else
      parameter load_delay = 300; // minimal load_unload time advance
   `endif

   initial begin

      //
      // --- establish a default time format for %t
      //
      $timeformat(-9,2," ns",18);

      //
      // --- default verbosity to 2 but also allow user override by
      //     using '+define+tmax_msg=N' on verilog compile line.
      //
      `ifdef tmax_msg
         verbose = `tmax_msg ;
      `else
         verbose = 2 ;
      `endif

      //
      // --- default pattern reporting interval to 5 but also allow user
      //     override by using '+define+tmax_rpt=N' on verilog compile line.
      //
      `ifdef tmax_rpt
         report_interval = `tmax_rpt ;
      `else
         report_interval = 5 ;
      `endif

      //
      // --- support generating Extened VCD output by using
      //     '+define+tmax_vcde' on verilog compile line.
      //
      `ifdef tmax_vcde
         // extended VCD, see IEEE Verilog P1364.1-1999 Draft 2
         if (verbose >= 2) $display("// %t : opening Extended VCD output file", $time);
         $dumpports( dut, "sim_vcde.out");
      `endif

      //
      // --- IDDQ PLI initialization
      //     User may activite by using '+define+tmax_iddq' on verilog compile line.
      //     Or by defining `tmax_iddq in this file.
      //
      `ifdef tmax_iddq
         if (verbose >= 3) $display("// %t : Initializing IDDQ PLI", $time);
         $ssi_iddq("dut AAA_tmax_testbench_1_16.dut");
         $ssi_iddq("verb on");
         $ssi_iddq("cycle 0");
         //
         // --- User may select one of the following two methods for fault seeding:
         //     #1 faults seeded by PLI (default)
         //     #2 faults supplied in a file
         //     Comment out the unused lines as needed (precede with '//').
         //     Replace the 'FAULTLIST_FILE' string with the actual file pathname.
         //
         $ssi_iddq("seed SA AAA_tmax_testbench_1_16.dut");   // no file, faults seeded by PLI
         //
         // $ssi_iddq("scope AAA_tmax_testbench_1_16.dut");   // set scope for faults from a file
         // $ssi_iddq("read_tmax FAULTLIST_FILE"); // read faults from a file
         //
      `endif

      POnames[0] = "hready_resp";
      POnames[1] = "hresp[1]";
      POnames[2] = "hresp[0]";
      POnames[3] = "hrdata[31]";
      POnames[4] = "hrdata[30]";
      POnames[5] = "hrdata[29]";
      POnames[6] = "hrdata[28]";
      POnames[7] = "hrdata[27]";
      POnames[8] = "hrdata[26]";
      POnames[9] = "hrdata[25]";
      POnames[10] = "hrdata[24]";
      POnames[11] = "hrdata[23]";
      POnames[12] = "hrdata[22]";
      POnames[13] = "hrdata[21]";
      POnames[14] = "hrdata[20]";
      POnames[15] = "hrdata[19]";
      POnames[16] = "hrdata[18]";
      POnames[17] = "hrdata[17]";
      POnames[18] = "hrdata[16]";
      POnames[19] = "hrdata[15]";
      POnames[20] = "hrdata[14]";
      POnames[21] = "hrdata[13]";
      POnames[22] = "hrdata[12]";
      POnames[23] = "hrdata[11]";
      POnames[24] = "hrdata[10]";
      POnames[25] = "hrdata[9]";
      POnames[26] = "hrdata[8]";
      POnames[27] = "hrdata[7]";
      POnames[28] = "hrdata[6]";
      POnames[29] = "hrdata[5]";
      POnames[30] = "hrdata[4]";
      POnames[31] = "hrdata[3]";
      POnames[32] = "hrdata[2]";
      POnames[33] = "hrdata[1]";
      POnames[34] = "hrdata[0]";
      POnames[35] = "so0";
      POnames[36] = "so1";
      POnames[37] = "so2";
      POnames[38] = "so3";
      CHAINnames[0] = "chain_1";
      CHAINnames[1] = "chain_2";
      CHAINnames[2] = "chain_3";
      CHAINnames[3] = "chain_4";
      CHAINpins[0] = "so0";
      CHAINpins[1] = "so1";
      CHAINpins[2] = "so2";
      CHAINpins[3] = "so3";
      SERIALM = 112'b0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
      INPINV[0] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      OUTINV[0] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      SHBEGM[0] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      INPINV[1] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      OUTINV[1] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      SHBEGM[1] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      INPINV[2] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      OUTINV[2] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      SHBEGM[2] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      INPINV[3] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      OUTINV[3] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      SHBEGM[3] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      nofails = 0; pattern = -1; lastpattern = 0;
      prev_pat = -2; error_banner = -2;

      if (verbose >=1) $display("// %t : Begin test_setup", $time);
      ->test_setup;
      #200; // 200


      /*** Scan test ***/

      if (verbose >= 1) $display("// %t : Begin patterns, first pattern = 0", $time);
pattern = 0; // 200
LOAD0 = 112'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
LOAD1 = 112'b0001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
LOAD2 = 112'b0001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
LOAD3 = 112'b0001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
UNLMSK[0] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
UNLMSK[1] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
UNLMSK[2] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
UNLMSK[3] = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
#0 ->load_unload;
#load_delay; // 500
ALLPIS = 62'b0110100011110100010111010000111100111001111100011111111011XXXX;
XPCT = 39'b100000000000000000000000000001001100000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture;
#200; // 700

pattern = 1; // 700
LOAD0 = 112'b0011101100100110100110100000101101001100001101011110101010101101111001111001101000000000001000000000000001000000;
LOAD1 = 112'b0100101010010100100010100000011111110110001101101111111111111011100111111101111111001111110011011101111111000001;
LOAD2 = 112'b0011101101100001010111001111010001010110111111111011010001011101011001000111110011100001010001011001101001010110;
LOAD3 = 112'b0010011101110011110100101111111000011011011110110101110000110101001111101011111001000111011101111011110100010010;
UNLOAD[0] = 112'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 1000
ALLPIS = 62'b01111111111111111111111111111111111100000001001111111111100001;
XPCT = 39'b100000000000000000000000000000000000100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 1300

pattern = 2; // 1300
LOAD0 = 112'b1001110010100011000111010101101000001100101010100110000110100011011110110111101111111111110111111111111111110110;
LOAD1 = 112'b0011000001110111100011101101101010100000011100111110011000110011111001111101000000101101110111100011110010111111;
LOAD2 = 112'b0010011110101101101111110001101110111000111000010101010000010000101010001101010110101101000000110000111011100100;
LOAD3 = 112'b0100111001111111110010011010000100101110011001101010101000001000001011010111011010110010001011100111011011111111;
UNLOAD[0] = 112'b0000001000100110100110100000101101001100101000000000001010001101101110000000001111111111111111111111111111111111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000001000000000000001000001101110111000000000001000000000000001000000000000000010000000000000010000010100000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000000100000000000000100000000000010000000000000010000000000001000001011100000000000100000000000000100000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000001101110000000000001000000000000100000000000000100000000000010000000000000010000000000001000000000000001000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 1600
ALLPIS = 62'b01110000000000000000000000000000000000000000110110000001100010;
XPCT = 39'b000000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 1900

pattern = 3; // 1900
LOAD0 = 112'b0101111001011100101000100000010111110011001110110110010100100001000101100110001111111111110111111111111110111111;
LOAD1 = 112'b0011011011000101110001100010010100111101010100001011011110001111101111100101001111001101111101110110111001111101;
LOAD2 = 112'b0000001101111000101001011011110010010101100000011000000001110111111101111100010011111010000101101011001011001000;
LOAD3 = 112'b0000010011010010110001010000001011111001111011010111010100001110111000100110110101011000011100010010100001110010;
UNLOAD[0] = 112'b1101110010101010011000011010001101111011001011001011001101011110110001000111110000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000001010111x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111111111111011111111111011111111111111101111111111101111111111111110111001000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100001111111111111110111111111111111011111111111011111111111111101111111111101111111111111110111111111110111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 2200
ALLPIS = 62'b01111111111111111111111111111111111100000011000100111111101011;
XPCT = 39'b000000000000000000000000000000000000000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 2500

pattern = 4; // 2500
LOAD0 = 112'b1101111110001011001101111111110100111111010110101111111111010100001100100000010000111010101001001011101101111111;
LOAD1 = 112'b0000001000001000100011001000111101011010101011101101000111100001100000101000011110110010011101001111110011000000;
LOAD2 = 112'b0111011101111101110001010101101001010010011011010011010001111100101011000001100000010101001100010001110000010100;
LOAD3 = 112'b0011110000000100010000000101001001110110001011001000111010101101110101010100101000100010111101111110111000011101;
UNLOAD[0] = 112'b1111111000111011011001010010000100010110100110100100111000110001001010110110010000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b111111110111111111111110111111110000001111111111110111111111111110111111111111111101111111111111101111110000110x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111111111011111111111111011111111111101111111111111101111111111110111100000011111111111011111111111111011111111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000011111111110111111111111011111111111111011111111111101111111111111101111111111110111111111111110111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 2800
ALLPIS = 62'b01111110001111000010000100011011100100000001000101100001101111;
XPCT = 39'b000100001111011001001110100111111001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 3100

pattern = 5; // 3100
LOAD0 = 112'b1001110001101011001001001000000010010110100011000001010100010011010010001001001100001100011100110101110010101110;
LOAD1 = 112'b0111110011001000101101010100000001010011010110010010111010011111011111010111100001001101100110111001011101000100;
LOAD2 = 112'b0111001100001000111001010001011011011111010000010001111001100111100011111010100100000110101000011111000001110111;
LOAD3 = 112'b0111111010101100001000000010100000111111000001100101001101110110101110110110011111001101110011001110100001101011;
UNLOAD[0] = 112'b0000000010000101001000111000000111010110001111111111110001001101100111010100101000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b001111011001001110100111111000001110000000000000000000000000000000000000000000000000000000000000000000001100000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010111010111110001110010100101011101011111000111001010010101110101111100001110101110110100011110000110000010100x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100000100011100101001010111010111110001110010100101011101011111000111001010010101110101111100011100101001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 3400
ALLPIS = 62'b01110111000111100001000010001101110000000000001100110001100111;
XPCT = 39'b000000000000000000000000000000000001111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 3700

pattern = 6; // 3700
LOAD0 = 112'b1011100010100100010011011100111010110100010000110010101011001010111101101000011111001100000000100011010100011110;
LOAD1 = 112'b0111100100110110010010011000000011110010000101001000010000000010000000111001101011010100011000000100100011100111;
LOAD2 = 112'b0100101100011110110101100101110100111010110100010111011101000011011011000111010011011011010101101110111010111111;
LOAD3 = 112'b0101010011110001001100111100001100111101010010010001100111110001101110010010111000000110011100101000000110100011;
UNLOAD[0] = 112'b0000011101101011001001001000000010010110011110010110110101011000110110101000000011100011110000100001000110111001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110000100110110011011100101110001101100000000000000000000000000000000000000000000000000000000000000000000001000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b101011101010111000011001110010101110101011100001100111001010111010101100010101011001001011101001111101111101011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000101010101110000110011100101011101010111000011001110010101110101011100001100111001010111010101110000110011100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 4000
ALLPIS = 62'b01111011011110110101010101001001110100000011001101100111101001;
XPCT = 39'b000000101001000010000000010000000111111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 4300

pattern = 7; // 4300
LOAD0 = 112'b0110000100000011001100101011001100011011001101111110110100011100100011001110101111100101000000000001101111001000;
LOAD1 = 112'b0101011101111110111001110111111011001001100011001101001100000101000010110110110101111010001100000110110010111000;
LOAD2 = 112'b0110010110001110001111101110010101000101111101011011110011001111110101111110101111111000111111111011010101001011;
LOAD3 = 112'b0000100101010101100110001110010010011110101100001001100011110000110111101001011100010011001111010100000011010001;
UNLOAD[0] = 112'b1011111110100100010011011100111010110100100100110111000101011000100001001000000000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110101101010001100000010010000010000000111110110011011101110110111010111111110111011110111111111110111100000011x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000110110001111110011000000000011011000111111001100000000001101100011100000000010100100001000000001000000011100x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000111100000011100110000000000110110001111110011000000000011011000111111001100000000001101100011111100110000000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 4600
ALLPIS = 62'b01101101101111011010101010100100111011111110011110110011100100;
XPCT = 39'b100000000000000000000000000000000000110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 4900

pattern = 8; // 4900
LOAD0 = 112'b1111111011101111101110110101101110111010111011101100001111111001000100100011101010111010101010101001011000100101;
LOAD1 = 112'b0010011001000011100100101111010001011011000111000111110010111111011100110111100101101101111011111010101101011101;
LOAD2 = 112'b0000010000000111011011010100100101110011001010001100001111000001010110110010101000101010100110000000000000100100;
LOAD3 = 112'b0001100100011001101011011010000001101101100001100111100001010010100110010011011100001111010100111101101001001100;
UNLOAD[0] = 112'b0110000000110111111011010001110010001100111001111111010011001000101001010110110000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001001000110110101110101001010101000101110110111001111000000100000001100100000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000011011100101111001100000000001101110010111100110000000000110111001010010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010101111011110011000000000011011100101111001100000000001101110010111100110000000000110111001011110011000000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 5200
ALLPIS = 62'b01110110001010101000100001011101010010000001000100100111100000;
XPCT = 39'b100000000000000000000000000101111111000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 5500

pattern = 9; // 5500
LOAD0 = 112'b1010000111100010100110100111101100111100000010000000000011100001001000010000101001011110010101100100101100010010;
LOAD1 = 112'b0011001110100001000000010100110001111100111000110111101001111100111111000000110010010101000000010000000011000001;
LOAD2 = 112'b0000001000000011100100100101011001110001111110011010001000000001000100001010001111000110000111000110101110101110;
LOAD3 = 112'b0011110100100100100101111101000000110010110100110010110000101001010111100001101110000111101010011110110100100110;
UNLOAD[0] = 112'b0000011100110100001111100110011111001110111111011100000011010111000101001000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010010100010010101110010101001001010001001010111001010100100101000100100010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100011001011100101010010010100010010101110010101001001010001001010111001010100100101000100101011100101010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 5800
ALLPIS = 62'b01110011000101010100010000101110101000000010000110010011101000;
XPCT = 39'b100111000110111101001111100111111001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 6100

pattern = 10; // 6100
LOAD0 = 112'b1111011100001110111111000011000110110111110000110001110000000011011111111101010100101101001010110010011010001010;
LOAD1 = 112'b0100110010111010010000000101000001001011111110111111111011000101101111110111000001101111100010100000001111000001;
LOAD2 = 112'b0000000100000001110010110111111000001000011001011010110101011111011011101000000011110000100001101001100011000001;
LOAD3 = 112'b0101010010010000000010111110110000010101011010011000011000110100101011010000110111000011110101001111011010010011;
UNLOAD[0] = 112'b1010000011100010100110100111101100111100011110000111011011000100101100010000001000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001010011000011011010100000000010011010100010101010001111100011001010010000000001x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001001010001000010111001010100100101000100001011100101010010010100010001110000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001010100100100101110010101001001010001000010111001010100100101000100001011100101010010010100010000101110010101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 6400
ALLPIS = 62'b01111001100010101010001000010111010100001000000111001001101100;
XPCT = 39'b000011100000110111110001010000000111101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 6700

pattern = 11; // 6700
LOAD0 = 112'b1101111011001100000010001111011111111101010010100110100101111011110010011010000111011100101111100000100110000101;
LOAD1 = 112'b0111111111111111011101011111011110001011011111111111101101111111110110111000110111110110111111010111010101100111;
LOAD2 = 112'b0011011001000001000101111100000011111100101110110001110100011100010111011111111111101110111111111111111111111111;
LOAD3 = 112'b0001110001110110110101010111100110100010111011111100001100001101111111111111101001101111001001010000000101101101;
UNLOAD[0] = 112'b0000011011000011000111000000001101111111010110110010101011001000011101000101100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100000110111110001010000000110001100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100100101000101001011100101010010010100010100101110010101001001010001000000011111011111111101100010110111111011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000110010010010111001010100100101000101001011100101010010010100010100101110010101001001010001010010111001010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 7000
ALLPIS = 62'b01111100001100010000110000000100100100000011100110011011101100;
XPCT = 39'b000100011011111011011111101011101011100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 7300

pattern = 12; // 7300
LOAD0 = 112'b1000010110000011100010000010111100010001111000100110010100111001100011110010101010100100011101111001110000000000;
LOAD1 = 112'b0001110010100101101011011011000100000010101000111100000001101100001010101010000110100000011101000010100111011010;
LOAD2 = 112'b0101100111110101110011010101010100011110101011100011110000111000000101011000010101111111010010111000111010100100;
LOAD3 = 112'b0010110000100011111100100100010010111000111001010100010110111110101111001100001101101101000110111000001000100100;
UNLOAD[0] = 112'b0000011101111010111001110101111100101111111111100000101011000010111100011000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000001011000011110111010111100000101100001111011101011110000010110000100011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100101110111101110101111000001011000011110111010111100000101100001111011101011110000010110000111101110101111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 7600
ALLPIS = 62'b01111110111011001101101100001101011100000011010100110011101100;
XPCT = 39'b000000000000000000000000000000000001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 7900

pattern = 13; // 7900
LOAD0 = 112'b0100010100111101001110011011110100000100011011010101010001000101011100010101011101010011001110011100111100000000;
LOAD1 = 112'b0000011100101001011010100110111100110001110110011110000110110111000101010100000011010000001110100001010001000101;
LOAD2 = 112'b0110100010011000111001101010101110001111010100110001111000011100001010100010000001011011110100111110001110101001;
LOAD3 = 112'b0101000111101100111110100010011001010100011101101010001011010111010111011000101110110000110101001001111000010001;
UNLOAD[0] = 112'b0000010010000011100010000010111100010001000000000101101001111110111000010110110000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100100011101111001110000000001001001000010100100011101111001110000000000101001000111011110011100000000010000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110011100000000101001001110111001110000000010100100111011100111000000010010101010010001110111100111000000000010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000101000101010010011101110011100000000101001001110111001110000000010100100111011100111000000001010010011101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 8200
ALLPIS = 62'b01111111011101100110110110000110101100000000000110011000100110;
XPCT = 39'b100110110011110000110110111000101010011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 8500

pattern = 14; // 8500
LOAD0 = 112'b1110001110000110111110101001000011110100101010010010001001001000000001110100100011100001101101000111111101000000;
LOAD1 = 112'b0100101100010010011111100000101011001010000000010010001010001101011100110001011110110011000001010011101011100000;
LOAD2 = 112'b0011110110111001001101011110001110100111011100100011010110111000000111111110110010000110101000111000000110011011;
LOAD3 = 112'b0000100100001011101010101110010110100001100010001011011011001101110100011101110011100000100110000000010010000000;
UNLOAD[0] = 112'b0000010001101101010101000100010101110001001100100010001000101101011010010101100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111001110000001010100100111011100111000000101010010011101110011100000000000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000010101001001110111001110000001010100100111011100111000000101010010011101110011100000010101001001110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 8800
ALLPIS = 62'b01111111010011110110101111001100011000000000000110110011101001;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 9100

pattern = 15; // 9100
LOAD0 = 112'b1010011100010010010111011100100000111011100111001001000011100000101100110100000001110000110110010011110110100011;
LOAD1 = 112'b0111001011000110000111111000001011110001000000001001000101000110101110011000101111011001100000101001110110011011;
LOAD2 = 112'b0001111011011100001110101111000011010011101111010001011011001100001001111111010100100100101010011110000001100010;
LOAD3 = 112'b0001010100110101111011011101000110110110111110101010001101010110001110001110111001110000010011000000001001000000;
UNLOAD[0] = 112'b0000000010101001001000100100100000000111001110011110111101011001110000110000111000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000010000011100001101101000111111101000000111000011011010001111111010000010011000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001111110100000111000110110100111111010000011100011011010011111101000010010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100101101110001101101001111110100000111000110110100111111010000011100011011010011111101000001110001101101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 9400
ALLPIS = 62'b01110111101001111011010111100110001100000000000011011001101100;
XPCT = 39'b100000000000000000000000000011101001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 9700

pattern = 16; // 9700
LOAD0 = 112'b0011010100000011010000001000101011101011010001001100010101011110010100011111101101110011010001100000011100010011;
LOAD1 = 112'b0011011001101001101000110111000101111011011010011001101000110101001001010111101000110111110110010111111010011001;
LOAD2 = 112'b0011110100111101011110111100110100001001000011010011110111000000000010011100011111011001011111000000000101101011;
LOAD3 = 112'b0010110010001100011001100010001000100011111111010110011101001110101101100100110111010010110000110001101110010000;
UNLOAD[0] = 112'b0000010110011100100100001110000010110011011111011100110101000001101110000000001000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001110100000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100111111010000011100011011010011111101000001110001101101001111110100000011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100110100111000110110100111111010000011100011011010011111101000001110001101101001111110100000111000110110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 10000
ALLPIS = 62'b01111011001001111000011111111100001000000101000100010011100100;
XPCT = 39'b000000000000000000000000000000000000000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 10300

pattern = 17; // 10300
LOAD0 = 112'b0001110011001011100001011010111010011010000000100110001010001010101011100111101111110011100010011001100101001000;
LOAD1 = 112'b0000011101000010010011000100111101101011110111010001111110001100111010110000001011000000111101001000111101000010;
LOAD2 = 112'b0101100100010110010110110101001011100100010110010110110001010010011011111100111101100110000010010111110100101011;
LOAD3 = 112'b0110111011100111000100101100111000110011001101001000011110100101111111011110001001100111111000111011010001011110;
UNLOAD[0] = 112'b0100110001000100110001010101111001010001111001010110101000011101101111110111111000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110011010001100000011100010011001111000000000000000000000000000000000000000000000000000000000000000000000000100x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000110001001011100101000100000011000100101110010100010000001100010010010110111001101000110000001110001001101x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000110110010111001010001000000110001001011100101000100000011000100101110010100010000001100010010111001010001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 10600
ALLPIS = 62'b01111101011001111001111011110001001000000001000101110111101000;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 10900

pattern = 18; // 10900
LOAD0 = 112'b0101100110001010000001001101100110001001101001100001100001000110001011011011011011111000110001101100110010100100;
LOAD1 = 112'b0110001101010010000110111001001110100100101110101001011111000110011111011100001101100000011110100101011101110101;
LOAD2 = 112'b0010010100001110110001111010110110101111100011011010010111110101111110100011111101111101110000110100100101011000;
LOAD3 = 112'b0101101001001111110010000110011000011101100011100100001111010010101111100111110010101010110111011110001111010011;
UNLOAD[0] = 112'b0000010000000010011000101000101010101110001110111001000100101001001101100111110110101100111100111101111000100101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110011100010011001100101001001000110000111110011100010011001100101001001111100111000100110011001010010010100000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110011010100101111100110001011001101010010111110011000101100110101001001011011111001110001001100110010100100111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111101011111001100010110011010100101111100110001011001101010010111110011000101100110101001011111001100010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 11200
ALLPIS = 62'b01111110101100111100111101111000100100000010000100111011100100;
XPCT = 39'b000000000000000000000000000000000000101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 11500

pattern = 19; // 11500
LOAD0 = 112'b1101100111001110111111011101100011100111011110010001011001100101110100101100011001111100011000010110011101010000;
LOAD1 = 112'b0000011011001001101101100111111001001000111101110100011111100011001110101100000010110000001111010010001110111111;
LOAD2 = 112'b0101001010000100000001001100100011110111001000100010101001111001001110101101101100100100101010010101000101000000;
LOAD3 = 112'b0000111110101010111001100011001000001110110100110011000111001001010111010011111001010101011011101111000111101001;
UNLOAD[0] = 112'b0101100010001010000001001101100110001001110111001010110101101011100011110111100111010110011110011110111100010010;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100100011000010111100010001100101100110110001100001000001000011001100101001000001x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011001101010010111110011000101100110101001011111001100010110011010100100111100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000110101001101111100110001011001101010010111110011000101100110101001011111001100010110011010100101111100110001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 11800
ALLPIS = 62'b01111111010110011110011110111100010000010010111100011101101010;
XPCT = 39'b100000000000000000000000000000000001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 12100

pattern = 20; // 12100
LOAD0 = 112'b0101111111110011011101010110111101111110101010011111011011110010110011111000110000111111001100001011000110101010;
LOAD1 = 112'b0101100111010110010001110101000110010001111100110010111111011110111111111101110011110111100110110111011101010000;
LOAD2 = 112'b0110100101000010011110111110110111111001110010000011110101000110011010101101100011000000001110101111001011001011;
LOAD3 = 112'b0001000110101011011100110001110000001011011110011000110011001100101011101001111100101010101101110111100011110100;
UNLOAD[0] = 112'b1101100001111001000101100110010111010010010000000101010011101001101010010000101111101011001111001111011110001000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000001011000000111101001000110001001000000000100000011010011100110000000111100011010100100000100011010001010011x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b101100110101000011111001100010110011010100001111100110001011001101010011001111110111010001111110001100111010110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000110000001100111110011000101100110101000011111001100010110011010100001111100110001011001101010000111110011000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 12400
ALLPIS = 62'b01110111101011001111001111011110001000100001001100001111101101;
XPCT = 39'b100000000000000000000000000000010110110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 12700

pattern = 21; // 12700
LOAD0 = 112'b1101011011111100101100110011011111001101001011000010011011011111110011001111011100011101100110100101100011010101;
LOAD1 = 112'b0111110110000101110000000100111011001100011111011101000111111000110011111011000000001100000011110100100001001111;
LOAD2 = 112'b0011010010100001110110011011011010001110010010101001000101011001001100010010110010001011011100110101100000101111;
LOAD3 = 112'b0001010111101001000001101011001111000001001100100010111011000010111001010100111110010101011110111011110001111010;
UNLOAD[0] = 112'b0000011010111101100110110101001111111001000011001000100110111001001001110101000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000101100000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010110011010100001111100110001011001101010000111110011000101100110101000001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000110101000011111001100010110011010100001111100110001011001101010000111110011000101100110101000011111001100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 13000
ALLPIS = 62'b01110011110101100111100111101111000101000001101110000111101110;
XPCT = 39'b100101100000000110000001111010010001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 13300

pattern = 22; // 13300
LOAD0 = 112'b1100111111110100000111100101010100010000100111010000111110101011000100110110011011000110111001101011010010101010;
LOAD1 = 112'b0001010110111011110101001000001110110100110101110011101001101010000111101110011111001101000111111001010010001011;
LOAD2 = 112'b0110110010010001000010100110111000100111111100101111111000001011100000111100110010110111100010111010101101111100;
LOAD3 = 112'b0010100101110011111011011110101011000110001111101110110101100101110101011101101101000100011000101010010000011001;
UNLOAD[0] = 112'b0000011000101100001001101101111111001100011010100001001001110001100000110111100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001011001101011000111110011000101100110101100011111001100010110011010100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000010001111100110001011001101011000111110011000101100110101100011111001100010110011010110001111100110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 13600
ALLPIS = 62'b01100001000111110110000111111000101100000011110100111101100101;
XPCT = 39'b100000000000000000000000000000000001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 13900

pattern = 23; // 13900
LOAD0 = 112'b1101011000110101011110000110000101100111100000011100011101001101110011110000011100101010010110011100000110010110;
LOAD1 = 112'b0110111110110110010110111011101001011101101000000110111010100011010101100111010010001101000101101110101000001011;
LOAD2 = 112'b0000000010101001010000111000000001110011001001101100010110110011010010101100111110111001101101001001001111101011;
LOAD3 = 112'b0100110011010001110010100010011111010111100110100101010100110011000100111001000100101100111111100010100000101000;
UNLOAD[0] = 112'b0000011010011101000011111010101100010011110101001001111000001110000110100110100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000110111001101011010010101011000110111000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010110101010100110001011100101011010101010011000101110010101101010101010011001100011011100110101101001010101011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000110010101100010111001010110101010100110001011100101011010101010011000101110010101101010101001100010111001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 14200
ALLPIS = 62'b01100000011110111110110111110011011000011010111111100000101000;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 14500

pattern = 24; // 14500
LOAD0 = 112'b1100111100000101111010101111101101001100000011001010111110100100110100100101001111011111000001000111101000001010;
LOAD1 = 112'b0111000100110111101100001111111101110000111010001111010101000111110000101101100111000101110100111100110100110111;
LOAD2 = 112'b0111011010000101110001110111011101011001010010001101000001101111101111110110111101111010011110110101110110011101;
LOAD3 = 112'b0001011100111110100111111001110011010111110110110111110000111000101111101011010000011000101100000110111000110000;
UNLOAD[0] = 112'b0000010110100101100101111010001011001110100100110100010101100001010110011000001000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001011001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111000011001011001010001011011100001100101100101000101101110000110010100000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111010110010100010110111000011001011001010001011011100001100101100101000101101110000110010110010100010110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 14800
ALLPIS = 62'b01111000110010011010101111110110100010010010011000001110101110;
XPCT = 39'b100000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 15100

pattern = 25; // 15100
LOAD0 = 112'b1001001100100010010011110100110000101110000100101010100101010000010001101001110111101101100000110011110000000110;
LOAD1 = 112'b0011110001001111011011100011110111101000011101000111101010100011111000010111110011100010111010010110011011010001;
LOAD2 = 112'b0011101101000010111000111011101111101100101010000110110000100111111011100111011111001111100111101101001101100111;
LOAD3 = 112'b0001001111110111110001111110111000111101010101111000010100110111010011110101101000001100010110000011011100011000;
UNLOAD[0] = 112'b0000011000001100101011111010010011010010111011011010011100111111111011010101010100011001001101010111111011010001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001111000000101110111100000100111100000010111011110000010011110000001001000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011101111000001001111000000101110111100000100111100000010111011110000010011110000001011101111000001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 15400
ALLPIS = 62'b01101100011001001101010111111011010001001001001100000111100111;
XPCT = 39'b100000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 15700

pattern = 26; // 15700
LOAD0 = 112'b0011101000001110101110011101000110100010011011110100010110101111010010000010000110111100111010100000010111000010;
LOAD1 = 112'b0000010111001001011111111001111000111111110100111110111111000101100010010000100110101010011011001100001111001001;
LOAD2 = 112'b0110101101100001000101101010010000100011000000101000001011110011010111101101010001100010101100011101110110101110;
LOAD3 = 112'b0000001010101100111001010110010111111001000010001011001000011101001011101101000110001000111000110110000110101000;
UNLOAD[0] = 112'b0000001000100010010011110100110000101110000001100000011000010000100010110110000110001100100110101011111101101001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100111100000011111011110000010011110000001111101111000001001111000000101011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111110111110111100000100111100000011111011110000010011110000001111101111000001001111000000111110111100000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 16000
ALLPIS = 62'b01111110110001100011011111110010100110111011100001111101100001;
XPCT = 39'b000000000000000000000000000000000000010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 16300

pattern = 27; // 16300
LOAD0 = 112'b1001111110100001101000000101000000100111001101101100001011010101101001001011001111011111011101000000001111100001;
LOAD1 = 112'b0101010100011111111110011000001011011111110010011000000000001000001011001010101010101010001010001010001000000000;
LOAD2 = 112'b0011010110110000100101011101011011000000001011111100001001011110000010010011111010111011110000101010101011101011;
LOAD3 = 112'b0001011011110001001100111011001011110100100100000101110100000110110001010110100011000100011100011011000011010100;
UNLOAD[0] = 112'b0000001000001110101110011101000110100010110110010100110110111010110000011000000111011000110001101111111001010011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000111001110111100111010100000010111000011101111001110101000000101110000110010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000111100001101111011101000000011110000110111101110100000001111000011001000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000000010011011110111010000000111100001101111011101000000011110000110111101110100000001111000011011110111010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 16600
ALLPIS = 62'b01101111011000110001101111111001010011011101110000111110101000;
XPCT = 39'b000000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 16900

pattern = 28; // 16900
LOAD0 = 112'b1101001001011111101111111110001111101100100010000010100000110001100000101101111010100100100100011001101000110001;
LOAD1 = 112'b0101101010000110100100110110101111100000100111010010100101100111100110111111110110110001100000110000000010011100;
LOAD2 = 112'b0110110000011001001010110110110000001101011110110101101010001001010101011110010101010010011111010111010110101101;
LOAD3 = 112'b0010100010111001111101110110010010100100110111100100010001000110111111111100100011101100111101111010001001001110;
UNLOAD[0] = 112'b0000011011110010001010100011011111010001011001100011001000101010001000000111010111101100011000110111111100101001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010101010101000101000101000100101011001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000011110001110111101110100000001111000111011110111010000000111100000011111001001100000000000100000101100101x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111110011101111011101000000011110001110111101110100000001111000111011110111010000000111100011101111011101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 17200
ALLPIS = 62'b01101111010001011101000011110011100111110001111111100001101110;
XPCT = 39'b000000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 17500

pattern = 29; // 17500
LOAD0 = 112'b1101101111000110001010111110010011000000001111100000100000110111010111000011001001010011010010001100110000011010;
LOAD1 = 112'b0011011010100011001001001101101010101001010011101001010010110011110011011111111011011000110000011000000011011101;
LOAD2 = 112'b0011011000001100101101011011010100000110101101011010110101010000101110101011000101010101100111100101110101101101;
LOAD3 = 112'b0110010010100100010101011101101111101010110011011001100011111101001100111110010001110110011110111101000100100111;
UNLOAD[0] = 112'b1100001010001000001010000011000110000010111011111010111100011001000011110110000000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100100100100011001101000110001001100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110011000011000101001010010011001100001100010100101001001100110000110010000101010010010010001100110100011000010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110111001010010100100110011000011000101001010010011001100001100010100101001001100110000110001010010100100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 17800
ALLPIS = 62'b01100111101000101110100001111001110011111000111111110000100111;
XPCT = 39'b000000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 18100

pattern = 30; // 18100
LOAD0 = 112'b1001111010110101111111101111111000111111110111011101111100110001000000010100100100101010101001100110010100001100;
LOAD1 = 112'b0010110110101010010010010011011100001101101001110100101001011001111001101111111101101100011000001100000011111011;
LOAD2 = 112'b0101101100000110010110101101100110000011010101101101001010111000010011010001100101010101011001111001011101011101;
LOAD3 = 112'b0100011011010010100100111100011110100000010010000101010100111100110001011111001000111011001111011110100010010011;
UNLOAD[0] = 112'b0110101011000110001010111110010011000000000101111110110111011011100000000111010000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b111101101100011000001100000000000000000001010011010010001100110000011010010100110100100011001100000110110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011001100001100010100101001001100110000110001010010100100110011000011010000001001110100101001011001111001101111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000000101001010010011001100001100010100101001001100110000110001010010100100110011000011000101001010010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 18400
ALLPIS = 62'b01100011110100010111010000111100111001111100011111111000101011;
XPCT = 39'b000000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 18700

pattern = 31; // 18700
LOAD0 = 112'b0000101100011110110111111101111101001111011110011111011110100001111110010111110010010110010100110011001110000100;
LOAD1 = 112'b0010101101101010100100100100111100000101110100111010010100101100111100110111111110110110001100000110000001100101;
LOAD2 = 112'b0110110110000010010011000100101010011011011000111110100000110100111100110101111001010101010110011110010111010111;
LOAD3 = 112'b0001101000001100110001011010011001001101100111000100100011010101010011101111100100011101100111101111010001001001;
UNLOAD[0] = 112'b0011011011011101110111110011000100000001011111110110010001010100101010010100110001111010001011101000011110011100;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b101010101001100110010100001101001010001100101010101001100110010100001101001010101010011001100101000011011010100x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001100110000111001010010100100110011000011100101001010010011001100001100001110010101010100110011001010000110100x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000011010010010100101001001100110000111001010010100100110011000011100101001010010011001100001110010100101001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 19000
ALLPIS = 62'b01110001111010001011101000011110011100111110001111111100100101;
XPCT = 39'b000000000000000000000000000000000000010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 19300

pattern = 32; // 19300
LOAD0 = 112'b1001000100000100110011110011100011001001000010001101111001101101100110110011011111111001010000100110000101111101;
LOAD1 = 112'b0000110110100010101001011100010011111101111100110101011011101100110110011001011111101100000000100011111011001001;
LOAD2 = 112'b0111110110001000010010111011011110111000001110010011010100010100000000001101110000000111011011111000000111100100;
LOAD3 = 112'b0010100000010000000010101011000110000010010011010101101111010111110111111001011010001100110001010001011000001011;
UNLOAD[0] = 112'b0000000001111001111101111010000111111001011111111100000100011011101111010000001000111101000101110100001111001111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100110011000010100101001010010011001100001010010100101001001100110000101001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100001101001010010100100110011000010100101001010010011001100001010010100101001001100110000101001010010100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 19600
ALLPIS = 62'b01101110000000001101001011001111100100100110011110100001100000;
XPCT = 39'b000000000000000000000000000000000001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 19900

pattern = 33; // 19900
LOAD0 = 112'b1001111100011000111111000100101100111110100001000010111100110111110011010000101011111110101000000011001010111101;
LOAD1 = 112'b0000001101101000001010010111000011001111010110111110101101110110110011101110100111011100000010110001110100001010;
LOAD2 = 112'b0111111011000101101110010100010100100100011000100011010101110110010010101010101000000100110110111110010001111011;
LOAD3 = 112'b0110110100000000000001000101110011000001001000101011100111101011111111111100101101000110011000101000101100000101;
UNLOAD[0] = 112'b1001000000000100110011110011100011001001111110011100011101111111001010010111100000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001111001111111001010000100110000101111101111110010100001001100001011111010000001x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001100010111111111110101000000110001011111111111010100000011000101111110001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010100110111111101010000001100010111111111110101000000110001011111111111010100000011000101111111111101010000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 20200
ALLPIS = 62'b01110111000000000110100101100111110010010011001111010000101000;
XPCT = 39'b100000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 20500

pattern = 34; // 20500
LOAD0 = 112'b0001100100111100000000001011011100011011110010101100100111110110011111011001111110000110000100000111100100100011;
LOAD1 = 112'b0110110101111000001011111001100110001011000011110010001101010111111011111111001000010111000000101011000100100011;
LOAD2 = 112'b0000001011101010111100011011100110010011011100110101110110101001011000000101100010000111010110000011100011111110;
LOAD3 = 112'b0101011001010001000010111001101011100010110010000001011100101010011000100111001100101111111101000101001110001001;
UNLOAD[0] = 112'b0000011000111010000101101111101101001111011111100110001011000000100000110100110000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001001001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000110001011110111111010100000011000101111011111101010000001100010111110010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100100101111110101000000110001011110111111010100000011000101111011111101010000001100010111101111110101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 20800
ALLPIS = 62'b01100101100000001110011001111100011101101111111001001001101100;
XPCT = 39'b000000000000000000000000000000000000101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 21100

pattern = 35; // 21100
LOAD0 = 112'b0111011101111010100000110111010101100110011011010111101010010110101001011010110000111000010010000101110111101101;
LOAD1 = 112'b0101111011111100001011101010000100101001111111000110111110101101000011101100111001101111000000010100111010100100;
LOAD2 = 112'b0011110011111100110110001001111101001110110001111110110001011011011101101001000100100111101110001001101011011010;
LOAD3 = 112'b0000101101011010100011100111110011111011001011010100000001000010111111001010111100011011001111110011111111001111;
UNLOAD[0] = 112'b0001100000111100000000001011011100011011110100100000010110011001011011000110000010110000000111001100111110001110;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100100001011100000010101100010100001000000010111010010110001010110011000101010011010011010111101011101001000011x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001111010010001100001000010000111101001000110000100001000011110100100001001100001111001000110101011111101111111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010101010011000010000100001111010010001100001000010000111101001000110000100001000011110100100011000010000100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 21400
ALLPIS = 62'b01101100110000001010000111110001101010010001100010000101101110;
XPCT = 39'b100000000000000000000000000000000000100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 21700

pattern = 36; // 21700
LOAD0 = 112'b1100101010011011100100100000001011111110101111101000001100100110110010010011010111100101011001100100110010001001;
LOAD1 = 112'b0111100000011101001011100100110010110000010010011111010101001111010011101010000010011111110000111000110110011100;
LOAD2 = 112'b0010001111110110101000100101000111000000000000000100100101000100101100100001000001001111100000001010001100010000;
LOAD3 = 112'b0000010001111000011011010000101011101010110111011110011011001010010101011100000100000001010110101000100111101100;
UNLOAD[0] = 112'b0000011000010101001001111011111110111010011111010101110101101001100000010111000110011000000101000011111000110101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b111000010010000101110111101101000101000000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001011111110110001110001001000101111111011000111000100100010111111101110001000011100001001000010111011110110000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100101011000011100010010001011111110110001110001001000101111111011000111000100100010111111101100011100010010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 22000
ALLPIS = 62'b01111000011000001000001000110111010001101110101111100011100111;
XPCT = 39'b000000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 22300

pattern = 37; // 22300
LOAD0 = 112'b0111000110101101011001000001000001100010011011101010100011010011000000001100010011110011101100010010011101000100;
LOAD1 = 112'b0001111000000101110010111001000101001001001001001111101010100111101001110101000001001111111000011100011001001011;
LOAD2 = 112'b0001000111111011010100001000101100100101100010010000110011001111010010110000111100010010111000010010100011000000;
LOAD3 = 112'b0010001011101011101001011100001101111111111010011111010111101111011100101110000010000000101011010100010011110110;
UNLOAD[0] = 112'b0010001010011011100100100000001011111110000110110001010110011110101010011000000000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001001101000101111001101100100100110100010111100110110010010011010001000000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011110011011001001001101000101111001101100100100110100010111100110110010010011010001011110011011001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 22600
ALLPIS = 62'b01111100001100000100000100011011101000110111010111110001100011;
XPCT = 39'b000000000000000000000000000000000000000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 22900

pattern = 38; // 22900
LOAD0 = 112'b0110110001000100011100101001010011000110001010010001010001110110110010000101111110000011100110001111000011011111;
LOAD1 = 112'b0000101000100011110101110010001010011001011000011010101110111111000010100011111111001011111100101101110111001101;
LOAD2 = 112'b0101101101010011001010111010000101011110010101100010001110100100100111011111110011000110110101111100101111010110;
LOAD3 = 112'b0110000011111100110110010101000100111101101110011010010100001000011101001100000110000110111101111111101110010111;
UNLOAD[0] = 112'b0000000001101110101010001101001100000000010110011000111101110111101001100100100110000110000010000010001101110101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110011101100010010011101000101000010000011110011101100010010011101000100111100111011000100100111010001010010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100100110100010111100110110010010011010001011110011011001001001101000100011001111001110110001001001110100010011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000011101001111001101100100100110100010111100110110010010011010001011110011011001001001101000101111001101100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 23200
ALLPIS = 62'b01100000000110001111001001000010010000111101110101011001101001;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 23500

pattern = 39; // 23500
LOAD0 = 112'b1001001000100101101000100100101110000101110100101000001001010011100101001001101111000010110011100111100001101101;
LOAD1 = 112'b0100001010001000011101011100101011000101101100001101010111011111100001010001111111100101111110010110111010111010;
LOAD2 = 112'b0011101010111011010100011111000110111111101101111011010111110001001011010011110000110100101101011111011011110011;
LOAD3 = 112'b0110111011111100001011101010100010010110110111001100011010000100001010110111001101100110010010011101101000111000;
UNLOAD[0] = 112'b0000010000101001000101000111011011001000111101100000110011000100100011100110000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000110000011100110001111000011011111100000111001100011110000110111110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011110001101111100000110011001111000110111110000011001100111100011011100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011000001100110011110001101111100000110011001111000110111110000011001100111100011011111000001100110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 23800
ALLPIS = 62'b01110000000011000111100100100001001000011110111010101100100100;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 24100

pattern = 40; // 24100
LOAD0 = 112'b0011101001010111110011011111100110100111001100110100111000111000011010010111111100011011001001010101111101001000;
LOAD1 = 112'b0111110100000010001110001011011110011010101010111011110000000011000110110001100000011110111111101000100101100000;
LOAD2 = 112'b0110000011010101000111000001001101101010001101001000110010001110001111100010000100001110010000101111110001011010;
LOAD3 = 112'b0100000011101110000111111110010011000101001001110010000010010101110110000010111100111111111000011111101100010111;
UNLOAD[0] = 112'b1011001000100101101000100100101110000101110110111111110101101001110010011000000000000001100011110010010000100100;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101000001000000000000000000000000000000000000000000000000000000000000000001010001x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001111000110111110000011001100111100011011111000001100110011110001101100011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000011111111100000110011001111000110111110000011001100111100011011111000001100110011110001101111100000110011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 24400
ALLPIS = 62'b01110110000001101110111001011111000000101001000011110111101010;
XPCT = 39'b000000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 24700

pattern = 41; // 24700
LOAD0 = 112'b0000101110111110100100011111100011101010111100010001101011100011101010001000101010001100100100111010110110100111;
LOAD1 = 112'b0101111101000010000011100010111001010000110101011101111000000001100011011000110000001111011111110100010010101111;
LOAD2 = 112'b0111000001101011010100010110111101001010010011101100001001001100100001000101011001000110100100011011101100010100;
LOAD3 = 112'b0000001010111010010011011111011001100010100001111000010001000010111111000001011010011111111100001111110110001011;
UNLOAD[0] = 112'b0000001000110011010011100011100001101001101110100100111010011111100110000100000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b011011001001010101111101001001000011000100011011001001010101111101001001000110110010010101011111010010010000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b101011110100101000110100100110101111010010100011010010011010111101001000000110001101100100101010111110100100100x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111101110001101001001101011110100101000110100100110101111010010100011010010011010111101001010001101001001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 25000
ALLPIS = 62'b01111011000000110111011100101111100000010100100001111011101101;
XPCT = 39'b000000000000000000000000000000000000110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 25300

pattern = 42; // 25300
LOAD0 = 112'b1111011011000101011110111001111110010101111110000100110101110000110101000001010101000111010010001101011111010000;
LOAD1 = 112'b0001011111010000100000111000101011100001110000001110011110001000011001001100011010101111101101010010000000010011;
LOAD2 = 112'b0111100000110101100101100111010111011110011110010110111111000000100101110111111110010100101001010110101111000101;
LOAD3 = 112'b0011101011100001010111100011100011111000010010101001001110100110001111100000101111001111111110000111111011000101;
UNLOAD[0] = 112'b0000001010111110100100011111100011101010011011100010111010101101001011000100110101100000011011101110010111110001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110101111010010100011010010011010111101001010001101001001101011110100101000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000000001000110100100110101111010010100011010010011010111101001010001101001001101011110100101000110100100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 25600
ALLPIS = 62'b01101101100000011011101110010111110000001010010000111101101110;
XPCT = 39'b000000000000000000000000000000000001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 25900

pattern = 43; // 25900
LOAD0 = 112'b0100100101010110101011101001000111010101011101011101100011010101111100010000011101011000111001000000100010010111;
LOAD1 = 112'b0010100001010110101001010010011000010001110001101010000101101100101110101111010011101111110111011110111100000011;
LOAD2 = 112'b0000000110010011001110100010011100010001010011010101111000001111100011100110010111100110010011101101111101010111;
LOAD3 = 112'b0110100111011110111110110100100010011110111111001011101011010011010100101001001101101011001110010010100101101001;
UNLOAD[0] = 112'b0000011001110111111010100010010000110010011000010101001011011110100111101000000110110000001101110111001011111001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011010111101001010001101001001101011110100101000110100100110101111010001011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111100010100011010010011010111101001010001101001001101011110100101000110100100110101111010010100011010010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 26200
ALLPIS = 62'b01101000110000000000111100000100011100100011010110111111101111;
XPCT = 39'b100000000000000000000000000000000000001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 26500

pattern = 44; // 26500
LOAD0 = 112'b1101101110000111011100111010001000100001101100101000000101110110110110101101010001010101001100110110010100110101;
LOAD1 = 112'b0110011110110111100011001000111001111001100100001000011001011010100001001110110110011011111011001100100100101000;
LOAD2 = 112'b0011110101000001010101110011000001001110111011110111001111110001011110010110101001111011111111100011011000110001;
LOAD3 = 112'b0101001000101001101101110010101000010100111100110000000000001000000110001101111100111001010110011000001010111111;
UNLOAD[0] = 112'b0100100001010110101011101001000111010101100010100001110000010100111100010100101000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000010100010011111010000011100110001100001101111101100001110101110011111100000011x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000001001001011010110011100100000100100101101011001110010000010010010100010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010111011110101100111001000001001001011010110011100100000100100101101011001110010000010010010110101100111001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 26800
ALLPIS = 62'b01111010011000001101010101001101101010110111110101111110100111;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 27100

pattern = 45; // 27100
LOAD0 = 112'b0001111011010010101110011111000001001000000110011111100100000011001100011000010000101011100110001011001110011001;
LOAD1 = 112'b0001100111000111010000111010000011101100111010001100001100101101011010100111010011101111110101001110011010100000;
LOAD2 = 112'b0101111010100001101010101010111101101111010010011011011011101101010011010101011110001011101110101101110111001011;
LOAD3 = 112'b0011101111100101011110010000101001100010100011011000001101010111010010000110111110011100101011001100000101011111;
UNLOAD[0] = 112'b0000001010110010100000010111011011011010001000110101110011110110111100010101100101001100000110101010100110110101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000001010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b101100110011010010101100110010110011001101001010110011001011001100110101010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000000101000101011001100101100110011010010101100110010110011001101001010110011001011001100110100101011001100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 27400
ALLPIS = 62'b01101101001100000110101010100110110101011011111010111111100011;
XPCT = 39'b100000000000000000000000000000000000010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 27700

pattern = 46; // 27700
LOAD0 = 112'b1101110001101011100001011110000011001010111100000100110110001110101110000111000111101101100011000011100110110010;
LOAD1 = 112'b0100001111011001011111010000111000010110000101111111011101111010011110001010110010001010111110010000110010000001;
LOAD2 = 112'b0111100101110110010101101111101100111101111010111110010100011111111001110011010011100100100100000010011010000101;
LOAD3 = 112'b0100101110001100101101100011000010111011000011111000101001011100001110001100100011000001010101010000110111010100;
UNLOAD[0] = 112'b0000011000101010000001101010000110111100101000100011010001001101101001001000000110100110000011010101010011011011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101101011000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010110011001100001010110011001011001100110000101011001100101100110011001001000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111100100010101100110010110011001100001010110011001011001100110000101011001100101100110011000010101100110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 28000
ALLPIS = 62'b01111000100110001110011110011100111110001011100011111110100001;
XPCT = 39'b100000000000000000000000000000000001111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 28300

pattern = 47; // 28300
LOAD0 = 112'b1111111010100101111000100111010000110100100000100011000101110111100000010010000111110101110001010001110011011000;
LOAD1 = 112'b0011000011110100110111110100001001010011000010110101000100010101100111100101011011001101110111100000110010100011;
LOAD2 = 112'b0000100101101100000010110111111010011110111110011111101010001011111100111011101100111000001001010000100110100001;
LOAD3 = 112'b0001001001110111010110110110101000001011000001011001010011001001111111011101000010100001010010011011101101010010;
UNLOAD[0] = 112'b0000010011110000010011011000111010111000001011010110001001000100111100110111010100010011000111001111001110011111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000010111000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000111011011001111011110001100011101101100111101111000110001110110110000011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000110001111110111100011000111011011001111011110001100011101101100111101111000110001110110110011110111100011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 28600
ALLPIS = 62'b01111100010011000111001111001110011111000101110001111111100000;
XPCT = 39'b000000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 28900

pattern = 48; // 28900
LOAD0 = 112'b0010110111000111010000011000001101001001010010000100011011010110010110110010101100000000101000111110110000010001;
LOAD1 = 112'b0010000110011111100100100001010011001000111101100010101100110010010001111011110011001110101111000111110100001001;
LOAD2 = 112'b0001111110011100100001101000101001100001001010101100111010111000011100001000010011001100011001111100011110001110;
LOAD3 = 112'b0010111110001111110001100011111010100100100001001011001101000000111110111101110110110110111111000101101111101000;
UNLOAD[0] = 112'b0000011001101000000000001110100101011001110111000001000000001000001001101000000110001001100011100111100111001111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001010100000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100011101101101111101111000110001110110110111110111100011000111011011000011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000101110111111011110001100011101101101111101111000110001110110110111110111100011000111011011011111011110001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 29200
ALLPIS = 62'b01100000001001101110101100101000101011000100100110011110100000;
XPCT = 39'b100000000000000000000000000000000000000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 29500

pattern = 49; // 29500
LOAD0 = 112'b0111010001001000000010100010000111011010001011011101110100000110101101101000000101111011000100101001011001110100;
LOAD1 = 112'b0100010111000101010000010100001110011101000010001100001101110101111110100100100110001011010111000000000010000001;
LOAD2 = 112'b0110001101011011010000000111001100011110110011110101100010110101101100000111111000110001011101100111010000000101;
LOAD3 = 112'b0100111001100001111010011010111011011000000011110001011001011111111000000010100101101110011001011000100010011010;
UNLOAD[0] = 112'b0000010011000111010000011000001101001001011000010011111100010011100001100000001000000100110111010110010100010101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101001000000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111101100001001000000010100011110110000100100000001010001111011000010010000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000010110010000000101000111101100001001000000010100011110110000100100000001010001111011000010010000000101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 29800
ALLPIS = 62'b01101110000100111010011101011011110001000100001101101110100000;
XPCT = 39'b000000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 30100

pattern = 50; // 30100
LOAD0 = 112'b1001111111001000100110000110101100010011110010100011101010000100101010110101001010111100100010100100101100111011;
LOAD1 = 112'b0011000101110001010100000101000111000111100001000110000110111010111111010010010011000101101011100000000010101111;
LOAD2 = 112'b0010000010001011001000000011101010001111011010111010110001011110110010001011100010001001010111001001110100000111;
LOAD3 = 112'b0001100011001010001000111001110001010101100010100101101101001110000000011001010011110001011110101111100111101101;
UNLOAD[0] = 112'b0000010001001000000010100010000111011010101000011100110011111011001010001000000111000010011101001110101101111001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b111011000100101001011001110101100011001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010010100111011011110100010001001010011101101111010001000100101001110101011110111101100010010100101100111010101x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000101100010111101000100010010100111011011110100010001001010011101101111010001000100101001110110111101000100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 30400
ALLPIS = 62'b01110111000010011101001110101101111000100010000110110111101000;
XPCT = 39'b000000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 30700

pattern = 51; // 30700
LOAD0 = 112'b1000101010001001000110100100001000000111100010111001011101000010101011010010001101011111010001000010011010011111;
LOAD1 = 112'b0110110001011100010101000001011000110111010000100011000011011101011111101001001001100010110101110000000010011110;
LOAD2 = 112'b0101000001000101011110110010001001010010101110001011101100101101111000001100100000100010010101100010011101000111;
LOAD3 = 112'b0010011101101000100110110110110010111010000110011100100110100111101110001100101001111000101111010111110011110110;
UNLOAD[0] = 112'b0000011111001010001110101000010010101011100010111011101111110111001111100101010000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001000001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001001010011100101111010001000100101001110010111101000100010010100111000011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100111001001011110100010001001010011100101111010001000100101001110010111101000100010010100111001011110100010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 31000
ALLPIS = 62'b01101011100001001110100111010110111100010001000011011011100100;
XPCT = 39'b100000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 31300

pattern = 52; // 31300
LOAD0 = 112'b0111000001110110001011100000001011110010010001011110101110100010010101100011101110101111101000110001000101001110;
LOAD1 = 112'b0111101100010101100101010000010111011111001000010001100001101110101111110100100100110001011010111000000000010010;
LOAD2 = 112'b0010100000100010001100101000110101101011110011001110010110000010001110000001011000001000100101001000110111010011;
LOAD3 = 112'b0111111011101001000011101011011101010101000110001111000011110011100111000110010100111100010111101011111001111011;
UNLOAD[0] = 112'b0111111110001001000110100100001000000111010111110000001100000110011000011000000101110000100111010011101011011110;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010010x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000100101001111010111101000100010010100111101011110100010001001010011111000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000000010101111010001000100101001111010111101000100010010100111101011110100010001001010011110101111010001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 31600
ALLPIS = 62'b01100101110000100111010011101011011110001000100001101101101010;
XPCT = 39'b000000000000000000000000000000000000101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 31900

pattern = 53; // 31900
LOAD0 = 112'b0001010010010011010000011001000101011001110110100001010101100001110001110110011111010101110100101000101010100101;
LOAD1 = 112'b0111111011000101011001010100001101110110100100001000110000110111010111111010010010011000101101011100000001101100;
LOAD2 = 112'b0100010010001111100111000000010110010001111001100111001010011010111011001000111010000010001001000010011101110000;
LOAD3 = 112'b0101100110101011100001010101111010101110100010000111110001011001110111001111011011111000001001111011111010111110;
UNLOAD[0] = 112'b0111000001110110001011100000001011110010101011110001101001100110001011001000000010111000010011101001110101101110;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010010011000101101011100000000101011001010100001011111111100001001100001000001110110110110100110001011000000010x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100010010100111101011110100010001001010011110101111010001000100101001100001000100001000110000110111010111111010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010111101011010111101000100010010100111101011110100010001001010011110101111010001000100101001111010111101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 32200
ALLPIS = 62'b01110010111000010011101001110101101111000100010000110110101101;
XPCT = 39'b100100100001000110000110111010111110111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 32500

pattern = 54; // 32500
LOAD0 = 112'b1111110010001011010110001111010001001011100011111000100110100100010100000100110100010010101010100010011100101111;
LOAD1 = 112'b0001001000010011111111001001011011000111101110111001000011110111011101100100010110100000010110001101111010111100;
LOAD2 = 112'b0100011100000110111011010011011011100110101001010000011010100000111111110010100010100111111001111000110000111110;
LOAD3 = 112'b0001010110110001110010010001101011011001000111010110010111111011001000110010000010110011010010000010111000001111;
UNLOAD[0] = 112'b0000011111011010000101010110000111000111010111001100010111101100111100110110100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001001111000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010001001010011110101111010001000100101001111010111101000100010010100100000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100110101011101011110100010001001010011110101111010001000100101001111010111101000100010010100111101011110100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 32800
ALLPIS = 62'b01100111011100000100111111110101010011000100010110111010101110;
XPCT = 39'b100000000000000000000000000100111111010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 33100

pattern = 55; // 33100
LOAD0 = 112'b1000111000000010010111011100001011001010100001011001110000101100010111000011100001110011000101000111001011101010;
LOAD1 = 112'b0100100100100100110110101110001110001010000001001001011010111111110000001001110100111100101011100111100101010011;
LOAD2 = 112'b0011011001001000010101011010110001011101000011001011000010101101110101101000101000101011100101100110011011101111;
LOAD3 = 112'b0001001111010100100110100111111010111101000100110010111100110101001010000101000101101101001011000100101011000001;
UNLOAD[0] = 112'b0000011110001111100010011010010001010000110000000011000110101111011001010101000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b001011010000001011000110111100000000001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000100110010111000100010101000010011001011100010001010100001001100101100000010111011100100001111011101110110010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000010001000101010000100110010111000100010101000010011001011100010001010100001001100101110001000101010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 33400
ALLPIS = 62'b01101101101110001111010100110101001101000100010101111100101111;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 33700

pattern = 56; // 33700
LOAD0 = 112'b1001011110010011110111111111100010011010110010101011000001111000101101011001001011000001110010010101100100001010;
LOAD1 = 112'b0111111111101001100100110111111010101101001001100101101110100111011010101110010111111010000111111011110011000111;
LOAD2 = 112'b0010011010101100100010011110000000000000110101000110111110101111011100111100110010001101100010110001110001011111;
LOAD3 = 112'b0010111100001011110011011111100010111000110100101011010101100000101001011011111000111010010100110011001101101011;
UNLOAD[0] = 112'b0000011001011110111001001111010001000110100111001101001110101010001001011000000110110111000111101010011010100111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001110001110100011100100010100111000111010001110010001010011100011101000000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111010100111001000101001110001110100011100100010100111000111010001110010001010011100011101000111001000101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 34000
ALLPIS = 62'b01111000110111001010100001010101000010000100010100011111101111;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 34300

pattern = 57; // 34300
LOAD0 = 112'b1110111001011000111101111111110100010101111001001011100000111110010110100001010101100000111001001010110010000101;
LOAD1 = 112'b0111111111111010011001001101110110001111001100101100011011110001000111100100111010010011100010100010000100011011;
LOAD2 = 112'b0101001101010110010001001111000000000000011001100001001111010111101110011011011100100010011000111100001100010111;
LOAD3 = 112'b0101010000100101100111101001011101110110101011110000011110101000010110001101111100011101001010011001100110110101;
UNLOAD[0] = 112'b0000011010110100101111011110101001101111011110011101011110001001110100000101010100011011100101010000101010100001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101110001011000001110010010101100100001010110000011100100101011001000010110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b101011010000100110000111001010101101000010011000011100101010110100001011000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100101101100001110010101011010000100110000111001010101101000010011000011100101010110100001001100001110010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 34600
ALLPIS = 62'b01101100011011100101010000101010100001000010001010001111101111;
XPCT = 39'b000000000000000000000000000011111011111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 34900

pattern = 58; // 34900
LOAD0 = 112'b1001010100111010101100110110001101101101111100101000111110100011001110011100001101001011001100110011010000111101;
LOAD1 = 112'b0111001001011110000111001111000110101011001110101110000010000101000000111010010010110000100001110111101101100100;
LOAD2 = 112'b0001000010001001000000010100110100101110011001010010011000000010010001011111001111001011111101110111000100100101;
LOAD3 = 112'b0001011111000101111111110101110100110100000011101110100010100011001100101110110111001010100001011001000001011010;
UNLOAD[0] = 112'b0000011001100110100001010101100001111011101000111100100110110000100111101000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000001001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010101101000011011000011100101010110100001101100001110010101011010000100011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100100110110000111001010101101000011011000011100101010110100001101100001110010101011010000110110000111001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 35200
ALLPIS = 62'b01111000001101111111100011011010110100000111011011100110101111;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 35500

pattern = 59; // 35500
LOAD0 = 112'b0111111001001101011010011011010011101110100010100001001100110100100110111111111010100100100110101001101100011100;
LOAD1 = 112'b0011110010010101100001110011111110011100100111010111000001000010100000011101001001011000010000111011110110011110;
LOAD2 = 112'b0100101000010000011100011000100100110011010101000100010110010110001000010100100011110110111111001101110001001101;
LOAD3 = 112'b0011110101011100101111111010111110010110000000110111010001110001100010011111110010000001001010001110110101101000;
UNLOAD[0] = 112'b0000011111110010100011111010001100111001101100101001100100111100111111110100010100000110111111110001101101011011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b001001011000010000111011110110100000000000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100110100011111010010100110010011010001111101001010011001001101000111101000000111010111000001000010100000011101x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000010100101001100100110100011111010010100110010011010001111101001010011001001101000111110100101001100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 35800
ALLPIS = 62'b01111100000110111111110001101101011010000011101101110011100111;
XPCT = 39'b100000000000000000000000000110011110010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 36100

pattern = 60; // 36100
LOAD0 = 112'b1000111111110000011101001110011011010000101011001100110111000000010111001100000110101010000011100010111111110011;
LOAD1 = 112'b0010001010000101110001000000100101111110001111010110111011001101100110010111111011000000001000111110000011010111;
LOAD2 = 112'b0101100010000000001100110110011011100101110000110111011001101001000000010100111100111110110100001011011011110011;
LOAD3 = 112'b0111001100101110000111110010101000101010100010111110111010001110000100010110100011001100010100010110000010111111;
UNLOAD[0] = 112'b0000011010001010000100110011010010011011101110000101100110100001101100110100000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010011010001110101001010011001001101000111010100101001100100110100011100000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100101011101010010100110010011010001110101001010011001001101000111010100101001100100110100011101010010100110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 36400
ALLPIS = 62'b01100000000011010010110011111001001001100111101000011000100011;
XPCT = 39'b100000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 36700

pattern = 61; // 36700
LOAD0 = 112'b0101010111111100000110110101011001110001000000010111110101000000001001100100110111010100000001110001011111111010;
LOAD1 = 112'b0110100010100001011100010000000011111011100111101011011101100110110011001011111101100000000100011111000001110111;
LOAD2 = 112'b0100011001000100000110011011000101110010111010011011011100100100101000010010010111001011101101010010100110111110;
LOAD3 = 112'b0111001110110100010010011011001000101010101100100111111011001111100001011111110100111001111000101100001001000110;
UNLOAD[0] = 112'b0000011110101100110011011100000001011100101111100011010110010100101000100100010000000001101001011001111100100101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000101111111001101010000001100010111111100110101000000110001011111110001000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011010100000011000101111111001101010000001100010111111100110101000000110001011111110011010100000011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 37000
ALLPIS = 62'b01110000000001101001011001111100100100110011110100001100100001;
XPCT = 39'b100000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 37300

pattern = 62; // 37300
LOAD0 = 112'b1010110101110010110110001110010101010111001001011011100110111110011011010011100111101001000000011000101111111110;
LOAD1 = 112'b0101101000101010010111000100101001111100110011110101101110110011011001100101111110110000000010001111100011111011;
LOAD2 = 112'b0111111101101000100011001101100010111001011100001101111110000110010000010110010001110010111011000100111001101001;
LOAD3 = 112'b0101000110010101001001001101100000011001010111010010111101101111100100100100100101010000100001000000011100101111;
UNLOAD[0] = 112'b0000011100000001011111010100000000100110101000111111111011010110010011010101000000000000110100101100111110010011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100010111111101110101000000110001011111110111010100000011000101111111000000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011101010000001100010111111101110101000000110001011111110111010100000011000101111111011101010000001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 37600
ALLPIS = 62'b01111000000000110100101100111110010010011001111010000110100000;
XPCT = 39'b100000000000000000000000000011101011111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 37900

pattern = 63; // 37900
LOAD0 = 112'b1110011010001111101000100111001101101100010111000010010100001100001111000101000111110110100000001100010011111111;
LOAD1 = 112'b0011011010001010100101110001001011101011111001111010110111011001101100110010111111011000000001000111110011100010;
LOAD2 = 112'b0111101100010001010101001100001000010110001011111000100011011101010011000111000000011101101110100001011110011000;
LOAD3 = 112'b0000101100010100100100010110100100000100101110101001011110111111100110110010110100011001100010000010110000010111;
UNLOAD[0] = 112'b0000010001110010110110001110010101010111011010111010101000001010101010000000001000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001010011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110001011111111111010100000011000101111111111101010000001100010111111100010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000110010111110101000000110001011111111111010100000011000101111111111101010000001100010111111111110101000000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 38200
ALLPIS = 62'b01111100000000011010010110011111001001001100111101000011100000;
XPCT = 39'b100000000000000000000000000000000001010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 38500

pattern = 64; // 38500
LOAD0 = 112'b1101101000100000110100110010001001000000111101001011111111100001000100001010100110000011111010000000001000110010;
LOAD1 = 112'b0011011001001111111001100011000110111100100001010111101100000110101101000011110110100101100110111110010100100101;
LOAD2 = 112'b0001101000111110100011111101110011011001010100110010011110011010111011010100000010111001101110100011101011101101;
LOAD3 = 112'b0100110100000111011010010111101001100011011100011100100101110000000000001101011001011110100111101001010111111010;
UNLOAD[0] = 112'b0000011001011100001001010000110000111100001100000110000110011101000010110101010110000000001101001011001111100101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100110000111110110100000001100010011111111111101101000000011000100111111111000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011000101111111111101010000001100010111111111110101000000110001011111101011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100010111111010100000011000101111111111101010000001100010111111111110101000000110001011111111111010100000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 38800
ALLPIS = 62'b01110011010101110001001110101000001111111000100100101100100000;
XPCT = 39'b100000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 39100

pattern = 65; // 39100
LOAD0 = 112'b1111111101011101111110110111111111111111111110110011111111110000100010001010000111000000111101100000000000011010;
LOAD1 = 112'b0000111100010001010100111010010111001010011000101001111110101010011100100011111001010000110011111111000000111100;
LOAD2 = 112'b0000110100011110010101111001110111011110001100100011011011110001110100101100000100111010001011111001101110101000;
LOAD3 = 112'b0000001000010101101110010110100000011000101010011101010010001101011000000110101100101111010011110100101011111101;
UNLOAD[0] = 112'b0000001000100000110100110010001001000000101010111010011100000010011010001000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000011111010000000001000110011000111011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000000011001100000111101000000000001100110000011110100000000000110000010111000001111101000000000100011001110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000111000001111010000000000011001100000111101000000000001100110000011110100000000000110011000001111010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 39400
ALLPIS = 62'b01101001101010111000100111010100000111111100010010010110100000;
XPCT = 39'b000000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 39700

pattern = 66; // 39700
LOAD0 = 112'b1001000011010000001010000100000000000000001111000010000100011001101000111101110001100001100100010000000000111111;
LOAD1 = 112'b0001110100101001100110000101000100001100011001000010010111000101100110010011001011001100111111010001110001111001;
LOAD2 = 112'b0101110010110001100010100100011011100010011000101100011110010100010000110000011110110111011000011001110001000100;
LOAD3 = 112'b0101100101010110111010100110001100100101000011110101101100011100111000101110001111001001001110010011000010000100;
UNLOAD[0] = 112'b0110111101100010000100001101011001001010000110101101000000001010001100110110010100110101011100010011101010000010;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000111101100000000000011011100000000000000000000000000000000000000000000000000000000000000000000000001010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000000001101110000011110100000000000110111000001111010000000000011011000011100000011110110000000000001101111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000000011100000111101000000000001101110000011110100000000000110111000001111010000000000011011100000111101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 40000
ALLPIS = 62'b01100111100000101101011101000010001100000110101101100111100000;
XPCT = 39'b100000000000000000000000000001100101011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 40300

pattern = 67; // 40300
LOAD0 = 112'b1010011111000011111110011111101111111111010110100010010111001100110110001101111010110001001000001000001000101110;
LOAD1 = 112'b0011000100000111000000000010010110111110001101110110100111100110011110001010010011000011111001010110101101000011;
LOAD2 = 112'b0011010001100110111110011100100001101110110110111101011010110111110101111010000001010000011000110101100111111000;
LOAD3 = 112'b0110010001011000011110101001110110011010101110010110100101001100000010111010011110111010000000100000110110111000;
UNLOAD[0] = 112'b0000000000111100001000010001100110100011110101100110100111001001100110010110000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100000000011110011000110010010000000001111001100011001001000000000111100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000101010100110001100100100000000011110011000110010010000000001111001100011001001000000000111100110001100100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 40600
ALLPIS = 62'b01100000100101100111100000001001001001111011110010011111100000;
XPCT = 39'b000000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 40900

pattern = 68; // 40900
LOAD0 = 112'b1100101111001011000010001000001000000000001100111010011100011111110110000101111011011011011110000100001000100100;
LOAD1 = 112'b0011101000001100101001100011100011100110000111101100111111110111100010000110111111000100011010010101000010001000;
LOAD2 = 112'b0000000000001101110100110011101011101110001101101100100011010101001101110100011010101100101000101110100010010001;
LOAD3 = 112'b0000000101101010001111000101011000011110011101110111000010110101000000110000010110000011100111111001001100100110;
UNLOAD[0] = 112'b0000011001011010001001011100110011011000001101101010111000100001001000010110001000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110001001000001000001000101111000111011010110001001000001000001000101110101100010010000010000010001011110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010000000010110101100100100001000000001011010110010010000100000000101110000101011000100100000100000100010111010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000101011001011001001000010000000010110101100100100001000000001011010110010010000100000000101101011001001000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 41200
ALLPIS = 62'b01100011000111000010111110101100101011000101011101100011101000;
XPCT = 39'b100000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 41500

pattern = 69; // 41500
LOAD0 = 112'b1011011000110001101001000100000001000000000001100110010000001011011001100001010001101110101111100010000000010011;
LOAD1 = 112'b0010111010000001101010011000110010111011000001110110011111010001011011100011011111001000001111101000100000001011;
LOAD2 = 112'b0000000000000110011010011001111001110111000111110110000001111010100010100010010110101010001010011011101000100000;
LOAD3 = 112'b0000101010101111101110001110011011110010010111011010011011111011000001011000001011000001110011111100100110010011;
UNLOAD[0] = 112'b0000001000110011101001110001111111011000100101111101001000011101011100000110000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001000000010010110110101111000100000001001011011010111100010000000100100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000101101001101101011110001000000010010110110101111000100000001001011011010111100010000000100101101101011110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 41800
ALLPIS = 62'b01110001100011100001011111010110010101100010101110110001101100;
XPCT = 39'b000000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 42100

pattern = 70; // 42100
LOAD0 = 112'b0100010011111011110100101011100111001111111101100000110111100101101000111001001010110100101101110001000000111010;
LOAD1 = 112'b0011110111101111100011000101001111100000000000101100100011111001010101100010011001010100100000011011000110101111;
LOAD2 = 112'b0101100011111001000110110001001111100010110111001001111110110111100010011110001111010011001100000101000001100001;
LOAD3 = 112'b0111110110110111100110100111111000111110011100010100001100101011000000110010101000111011001111100010111001100110;
UNLOAD[0] = 112'b0000011010100100010110101110100001011011010100000001111100010011010001001000000000110001110000101111101011001011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100111000000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000100000001000011011010111100010000000100001101101011110001000000010000010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000010101100110110101111000100000001000011011010111100010000000100001101101011110001000000010000110110101111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 42400
ALLPIS = 62'b01101011100100000001100001000011000101001001110011110100101110;
XPCT = 39'b100000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 42700

pattern = 71; // 42700
LOAD0 = 112'b1010011001000110101011111111110111110111111110111001011011110011110100011011110101011011010110011000101000011101;
LOAD1 = 112'b0010111101111001111000110001011110101001101000011110010011011110000010010011000110101000010000100111100010111111;
LOAD2 = 112'b0110110100011110001011011000100011110001011011100100111111011111010001001101000011110101110011000001000000011100;
LOAD3 = 112'b0100010110010101110010100011001010101101000000110010100000010010010110100000101110011111001111001011100010011001;
UNLOAD[0] = 112'b0000010011111011110100101011100111001111111011000001011111111111101011111000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100010000011100101101010110110001000001110010110101011011000100000111000010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100110110101011010101101100010000011100101101010110110001000001110010110101011011000100000111001011010101101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 43000
ALLPIS = 62'b01100101110010000000110000100001100010100100111001111010101111;
XPCT = 39'b100000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 43300

pattern = 72; // 43300
LOAD0 = 112'b1010010101001110011001010010101110100000000010010101010010011011111110001011010100101101010001101100011000111101;
LOAD1 = 112'b0011110110010001000111101111011000110001000001011100100100111010111000011011010000110000101110111000100101011011;
LOAD2 = 112'b0000000101110011100110010001100010100001111000000000110001100001000111100001111010000000110010010011111011101000;
LOAD3 = 112'b0110000100010101010100111100110110101110110001011111010110011000100100100011101010110101010111110100001111110100;
UNLOAD[0] = 112'b0111011000100111101100111010110001000100111101000010101010101000011111001000000000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b011011010110011000101000011101000000000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110001000001111010110101011011000100000111101011010101101100010000011110000010101101101011001100010100001110101x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000010101101010110110001000001111010110101011011000100000111101011010101101100010000011110101101010110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 43600
ALLPIS = 62'b01100001101100110001010110111000111110101010111000010001100111;
XPCT = 39'b100000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 43900

pattern = 73; // 43900
LOAD0 = 112'b1110011111101001010001011010000000100010000001000100101001001100111111001010101010010111101000010110001100011110;
LOAD1 = 112'b0000111101100110010001111011110001001100101010101100010000110111011110000101101010011000110101011100011001100010;
LOAD2 = 112'b0011011001011001001111010000100001001000001101000000011100001010101110010011101010100000001100100100101110111110;
LOAD3 = 112'b0110100000010010101010001110011111010011011100101110111011000100010110111110100111001000100000000110010011011011;
UNLOAD[0] = 112'b1111010001001110011001010010101110100000111000010111000010000001100000100000001000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000110100100101101010001101100011000111101001011010100011011000110001111010000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011000100011111001011101000101100010001111100101110100010110001000111100001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100010110010111010001011000100011111001011101000101100010001111100101110100010110001000111110010111010001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 44200
ALLPIS = 62'b01100000110110011000101011011100011111010101011100001000100011;
XPCT = 39'b000000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 44500

pattern = 74; // 44500
LOAD0 = 112'b0101001101110101100100100111000000001000110011001111010101110110000010000101101101001001110100101011000010001111;
LOAD1 = 112'b0100001111011011000100011110110000100010100000010111001001001110101110000110110100001100001011101110001010100011;
LOAD2 = 112'b0101101100101100000101111110001001111110111101110000000001101001010110111100111110101100000011001001001011101011;
LOAD3 = 112'b0100100000000110010101100111001011101101101011010110011101101010001011111111010011100100010000000011001001101101;
UNLOAD[0] = 112'b0000011011100011000011010011100110010101000110110011010011100111000111100110110000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000010011010010111101000010110001100011110100101111010000101100011000111110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b101100010001110100101110100010110001000111010010111010001011000100011100011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100010001001011101000101100010001110100101110100010110001000111010010111010001011000100011101001011101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 44800
ALLPIS = 62'b01100000011011001100010101101110001111101010101110000100101001;
XPCT = 39'b000000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 45100

pattern = 75; // 45100
LOAD0 = 112'b0101111110010101001101000110001111111011010011101111011000000011001101011110010000100111000000000101100001110111;
LOAD1 = 112'b0100011010111001001010100100100100100101110001011100001000100011111010000000101100100011100011101001010000000100;
LOAD2 = 112'b0111011110101001101000010100100110000000001110010010101010111110011010101010001101010111101110010001111001010011;
LOAD3 = 112'b0110000101010011000111011110111001011011100011010001011011000111010001010010110000101100101111101000110011001100;
UNLOAD[0] = 112'b0000001011001100111101010111011000001000110011110000100111010001110100010101110000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010110001000111010010111010001011000100011101001011101000101100010001110000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100101010100101110100010110001000111010010111010001011000100011101001011101000101100010001110100101110100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 45400
ALLPIS = 62'b01110011011000010111000100011111001000001101110011101110100100;
XPCT = 39'b100000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 45700

pattern = 76; // 45700
LOAD0 = 112'b1111011011100001011111101110101100000010010000100010011011100110000000001100000010010010011010100010111000001011;
LOAD1 = 112'b0100011111100011001011101010000110110010111001111001101000010101010000000011100000110100010111011010111110010011;
LOAD2 = 112'b0010000111101010000011011010000101111111111000011011110000010010000100110100010101101000010101010111100101111001;
LOAD3 = 112'b0010000100001111100010101000000000111111111001000110001010111101001010100100000001001000110000011101001110011100;
UNLOAD[0] = 112'b0000011001001110111101100000001100110101011000001101010010101101010011000110100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100111000000000101100001110111000000001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001011000111010001001100000000101100011101000100110000000010110001110110000000010011100000000010110000111011000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000000010011000000001011000111010001001100000000101100011101000100110000000010110001110100010011000000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 46000
ALLPIS = 62'b01101010111001111010101100100111101011111110011101011011100010;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 46300

pattern = 77; // 46300
LOAD0 = 112'b1111111011110100100111111101010111000000011111001101101100000010111000111111100101001000001101100001011100000110;
LOAD1 = 112'b0011000111111010010010111010100011011001011100111100110100001010101000000001110000011010001011101101011101001110;
LOAD2 = 112'b0001000011110101100101010100001110111010000000101101111011010001011010100010010001011110000101000101111001011100;
LOAD3 = 112'b0110000001110110110111101001000010000010010100001001110100100000111100010010000000100100011000001110100111001110;
UNLOAD[0] = 112'b0010111001000010001001101110011000000000110101000100001000110001001111010100010000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010010011010100010111000001011000110100000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000101100000100100100001101000010110000010010010000110100001011000001000010101001001001101010001011100000101010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100001101001000011010000101100000100100100001101000010110000010010010000110100001011000001001001000011010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 46600
ALLPIS = 62'b01110101011100111101010110010011110101111111001110101101100001;
XPCT = 39'b000000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 46900

pattern = 78; // 46900
LOAD0 = 112'b1001111001000101101100100001000101001111101111100000011110110110010000010000101000100101111100010000100110110000;
LOAD1 = 112'b0001100000010001010101000101000111011000000101101011111110000011010001101001101110100010101011100010110010011101;
LOAD2 = 112'b0001001001000101000101000000100000000100000100011001100011000000000011000110000011101110001111100011100101111101;
LOAD3 = 112'b0000011111011101000110111001111001100000011100111110101111101010011110100100011001001100101011101110000100011101;
UNLOAD[0] = 112'b0000011001111100110110110000001011100011011000100110100011101000011100010111110000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000101001000001101100001011100000111010010000011011000010111000001110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000010110000011010010000110100001011000001101001000011010000101100000100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000010100100001101000010110000011010010000110100001011000001101001000011010000101100000110100100001101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 47200
ALLPIS = 62'b01101001111011101111100101100001110101000111000011111010101000;
XPCT = 39'b100000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 47500

pattern = 79; // 47500
LOAD0 = 112'b1111111010100010110010011000100010100110001110100011000101111110111100100110100000010011111110001000010011011000;
LOAD1 = 112'b0000111010001110010111010011011111100001100111100100111011000000111100100001100111010100110001100100011111011101;
LOAD2 = 112'b0100100100100010000101100110100101001001110001110011000101000110100000000010010101101010100011111100111101011000;
LOAD3 = 112'b0001000001111000100011001100111100111000001011011110010111111101001011110010001100100110010101110111000010001110;
UNLOAD[0] = 112'b1100011001100000111110101101101101100001001001111101001100010111010010001000000100111101110111110010110000111010;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100101111100010000100110110001100000000000000000000000000000000000000000000000000000000000000000000000000010110x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100001011011000001001111110010000101101100000100111111001000010110110001000000010010111110001000010011011000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000000000010011111100100001011011000001001111110010000101101100000100111111001000010110110000010011111100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 47800
ALLPIS = 62'b01100100111101110111110010110000111010100011100001111101101100;
XPCT = 39'b000000000000000000000000000101111111010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 48100

pattern = 80; // 48100
LOAD0 = 112'b0001110011011011001011111010000010000111000110100101111000001101100000000001110110001001000101100100001101011111;
LOAD1 = 112'b0011010111101100011100010111110110010001110010100101110001100100110011010011000101001111101110001100011011111001;
LOAD2 = 112'b0110111000000101000001001111001001111000111101101111011110111010010001110111011011100111000110001100110100111101;
LOAD3 = 112'b0100111011101101011100111011000110111101010011010101011110000100100001000011110110000001100100010100000010101011;
UNLOAD[0] = 112'b0000011000111010001100010111111011110010000011001010101011101000101011010110110000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010000101101100000100111111001000010110110000010011111100100001011011000000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000000001001111110010000101101100000100111111001000010110110000010011111100100001011011000001001111110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 48400
ALLPIS = 62'b01110001001011001010110111110000010010101001010100010010100110;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 48700

pattern = 81; // 48700
LOAD0 = 112'b1100001010111100000101011001010010000101000000010000101010111011110101111101111001000101011000010010000010011100;
LOAD1 = 112'b0001101100110100011110100110111001111001111000000101010100110110110100101010010100000010010001111000011011001000;
LOAD2 = 112'b0100010101101001001011011010010011100101001011000101000001010111110111111010111100000001011111010000100110100100;
LOAD3 = 112'b0111011110111010000000100100001010111101101001111100111000011100101000010111010110111000010001000000001100100100;
UNLOAD[0] = 112'b0111110011011011001011111010000010000111010101011011010111101010011101001000000000100101100101011011111000001000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b001001000101100100001101011111100010100110001001000101100100001101011111100010010001011001000011010111111010101x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001000010101111100010100010100100001010111110001010001010010000101011101011011000100100010110010000110101111110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000011101111000101000101001000010101111100010100010100100001010111110001010001010010000101011111000101000101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 49000
ALLPIS = 62'b01101011110000010100010101010000000110101100001110100101101011;
XPCT = 39'b100000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 49300

pattern = 82; // 49300
LOAD0 = 112'b0011111101011111000000110110101000010010011111010101100001110001011010000011110000100011101100001001000001001101;
LOAD1 = 112'b0000111011001101100111101011101101101101011110001010100000111011010000110101001010101001001000110100001110100001;
LOAD2 = 112'b0010001010110101101010111011010101000001100100011011000100000011010100010011001010010001000111110100011000101011;
LOAD3 = 112'b0101110110100110111001110000001101111111111001001001100101100100011010101011101011011100001000100000000110010010;
UNLOAD[0] = 112'b0000001000000001000010101011101111010111001110011100001111011001100010100110000101111000001010001010101000000011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100100001001110010001101100010010000100111001000110110001001000010011100010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000010111000100011011000100100001001110010001101100010010000100111001000110110001001000010011100100011011000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 49600
ALLPIS = 62'b01100101111000001010001010101000000011010110000111010010100101;
XPCT = 39'b100000000000000000000000000000000000001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 49900

pattern = 83; // 49900
LOAD0 = 112'b1011111100101011101000001011010101000001101111100100110000011000101101001000111000010000110110100100100000100101;
LOAD1 = 112'b0110100100110011010011110010011100101111111110100001110101100111100111100010101101001010100110011100101110100101;
LOAD2 = 112'b0001000101011010001011111101000101110101011011001001000010111100101011011101100110100001000001101101010010001001;
LOAD3 = 112'b0010100111010110011100111000010010111111111101100100100010111010001001010101110101101110000100010000000011001001;
UNLOAD[0] = 112'b0000011010001110100100011010001100101111000110111110101010110010100110100000001000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100101010100100100011010000110001101001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010010000100110001000110110001001000010011000100011011000100100001001100011001111000101010000011101101000011010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000110100100010001101100010010000100110001000110110001001000010011000100011011000100100001001100010001101100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 50200
ALLPIS = 62'b01100010111100000101000101010100000001101011000011101001101010;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 50500

pattern = 84; // 50500
LOAD0 = 112'b1110010101000101111010000101101010100000100111100100000101111100010101011111001000001000011011000010011000010000;
LOAD1 = 112'b0001100001101110011100011110101010011111111111000000101010100110110110100101010010100000010010001111000000010110;
LOAD2 = 112'b0111100010111101100011011011010001011100100000101000010100001010110111101101111001111101000001001010010101100110;
LOAD3 = 112'b0110111001011111011110001100011001010111111111110010000001110101010000110001111111010011001111001001010000000101;
UNLOAD[0] = 112'b0000011100000101000001100100111111101001111101110011010110110010001010010000001000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010000110110100100100000100101000101001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001001000010010000100011011000100100001001000010001101100010010000100100001100001000011011010010010000010010000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100111011000001000110110001001000010010000100011011000100100001001000010001101100010010000100100001000110110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 50800
ALLPIS = 62'b01110001011110000010100010101010000000110101100001110100100101;
XPCT = 39'b000000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 51100

pattern = 85; // 51100
LOAD0 = 112'b0101011101100010110111000000110101011000001011101110001100001101001011010011010000000100001101010001000100001011;
LOAD1 = 112'b0100011000011001100111000111100111010110011101100010011111010001010001111000101011010010100011101111100001111010;
LOAD2 = 112'b0010010001010110111101001100111100111111001100101101101000000111001011111011100110011111010000010010110101011011;
LOAD3 = 112'b0101010000111010111111000110001000101111111011111001010000011010111000110101011101011011100001000100000000110010;
UNLOAD[0] = 112'b0100011110011110010000010111110001010101010011101001001100001110010101100111010000101111000001010001010101000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100011001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000100100001000000010001101100010010000100000001000110110001001000010011001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100101011100000100011011000100100001000000010001101100010010000100000001000110110001001000010000000100011011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 51400
ALLPIS = 62'b01101000101111000001010001010101000000011010110000111010101010;
XPCT = 39'b000000000000000000000000000010010100101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 51700

pattern = 86; // 51700
LOAD0 = 112'b1101010110011111100000101111110001011010001111110111011001001000011001101101011010000000111100011000101010110111;
LOAD1 = 112'b0100011111001001000000010010110011001110111110100111100110101101000000101010100010001101100010011101100111001011;
LOAD2 = 112'b0001111100100001100111001011001001001110011100111000011011011010011100110000110111011010011010110111000110111111;
LOAD3 = 112'b0110100011100010000010111110001000111010101001000111101101011111001100101110111101000000010000010011010110100000;
UNLOAD[0] = 112'b0000011011110100100000111101000001111011001111100011001010000011001100000111100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001101111000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100010010000100000001000110110001001000010000000100011011000100100001000011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100111000000010001101100010010000100000001000110110001001000010000000100011011000100100001000000010001101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 52000
ALLPIS = 62'b01110111000010010001100110000010101111110101111100110001100101;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 52300

pattern = 87; // 52300
LOAD0 = 112'b0001010000100110100000000110010011001011000001000011100011010000010100110011100011000001100100001100011001101001;
LOAD1 = 112'b0100011110111101001001100111101110001111011110000100011111010010001101010110100111100011010111110000100100001110;
LOAD2 = 112'b0110011111101100111000011000010011111110011011001110010011110011110101001110011111001010001000001110001010000010;
LOAD3 = 112'b0010010111001010001100000010011000111100000011011001110011110101100010010110101010011011001000011111011101110111;
UNLOAD[0] = 112'b0000010000111111011101100100100001100110011001110011100000010111001010100101100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000010011010000000111100011000101010110110100000001111000110001010101101110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110001001011010100000011110011000100101101010000001111001100010010110100000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111100001000000111100110001001011010100000011110011000100101101010000001111001100010010110101000000111100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 52600
ALLPIS = 62'b01111000110100111001111101101001011000000010011010110100100010;
XPCT = 39'b100000000000000000000000000000000000110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 52900

pattern = 88; // 52900
LOAD0 = 112'b1111111110011111111101101100111111001010011101101010001110001011001110000010100111100001001000000110001100000100;
LOAD1 = 112'b0100010100100010100011011010111000101010101100111101100001100111100011001000101101011110101101101110101110111000;
LOAD2 = 112'b0111010100100101101010110110111110100110000101010001111000101110101001110111000100011110001100100101011001001000;
LOAD3 = 112'b0010100100101101001011001100000000111111010010010111101100100000100101000110001000001101000001101111001001111111;
UNLOAD[0] = 112'b0000011100100110100000000110010011001011100101011100000100010101001011001000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000001100100001100011001101001000000001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011000100110100110000110010001100010011010011000011001000110001001101000000001100000110010000110001100110100011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000001100001100100011000100110100110000110010001100010011010011000011001000110001001101001100001100100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 53200
ALLPIS = 62'b01101111001111101101110000011100100011111001101001110110101001;
XPCT = 39'b100000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 53500

pattern = 89; // 53500
LOAD0 = 112'b0101001000000011111101101101110001011111100110101011000111000110100111001000100011110010100100000011000010000010;
LOAD1 = 112'b0011100111101010000010111110100010011001100111001010110001110110110101110100010010101010000110100011000011000010;
LOAD2 = 112'b0111101010010011010001110001111101001100110100111011001111101111001000011101101101010110110011001000000010010001;
LOAD3 = 112'b0100100010110111100101010110000000010111101100001011010110110000000110000011000100000110100000110111100100110111;
UNLOAD[0] = 112'b0001011010010001000001000001011000110010000110101001100110011011100001110110110000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000101000000000000000000000000000000000000000000000000000000000000000000000000100x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001100010000011111000100100000110001000001111100010010000011000100000100011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100101111110001001000001100010000011111000100100000110001000001111100010010000011000100000111110001001000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 53800
ALLPIS = 62'b01110111100111110110111000001110010001111100110100111011100100;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 54100

pattern = 90; // 54100
LOAD0 = 112'b1101001101100010000010000001100100000100010010000101100110010110001001011100010011111011101000100001101001110011;
LOAD1 = 112'b0001100000110111011001001100101101111001010010110010110100111111110111111001111111110000100101101111110100001101;
LOAD2 = 112'b0110011101110111110010000001101100110000110011110111110011110101000010011100110101101100000010010001111011001111;
LOAD3 = 112'b0100100110010011100000100110001100101010011001011110100101000100011010101100111011011101110111110010100101100101;
UNLOAD[0] = 112'b0000001000000011111101101101110001011111010110111111110001010011001011111000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000011000011110010100100000011000010000010111100101001000000110000100000110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000110001000000111100010010000011000100000011110001001000001100010000010001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100011001111000100100000110001000000111100010010000011000100000011110001001000001100010000001111000100100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 54400
ALLPIS = 62'b01111000100110001010010010101111000111000110111110110001100010;
XPCT = 39'b100000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 54700

pattern = 91; // 54700
LOAD0 = 112'b1001110001100100001001000000100110000010110001110011011110101100110111011111110101111110110100100000111000111011;
LOAD1 = 112'b0110011000001111010110010011001011101100101001011001011010011111111011111100111111111000010010110111111000110011;
LOAD2 = 112'b0011101110110101111001000000111010011000011010111011111001111110100001001011000101011110000000110100001110110111;
LOAD3 = 112'b0010010000000100110111111011010000011011010010111110011111110101000001101111000111100010110011000110100111000111;
UNLOAD[0] = 112'b0000000001001000010110011001011000100101111100011110101011010010101101110000101000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b111011101000100001101001110011001111000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000011000111000111110110100000001100011100011111011010000000110001110010011001111101110100010000110100111001011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110110101111101101000000011000111000111110110100000001100011100011111011010000000110001110001111101101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 55000
ALLPIS = 62'b01101100010011000101001001010111100011100011011111011000101001;
XPCT = 39'b000000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 55300

pattern = 92; // 55300
LOAD0 = 112'b1001001011011101111111111111111001101111101100101100100100111001101000101111110000111110100000100000010100101101;
LOAD1 = 112'b0100111111001110001100000111110010010110010101111011000001001011010000111101101001011001101111100101101011111101;
LOAD2 = 112'b0010001111100011011111011101101110010101011010101111100010100101100011100001110011101110001110111110101000000100;
LOAD3 = 112'b0010101100010110001011001100000000010011101101100011100100010010100101010110010111101001111010010101111110100011;
UNLOAD[0] = 112'b1110101111000111001101111010110011011101010010111101001100100110110100010000001000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001101011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000001100011101011111011010000000110001110101111101101000000011000111010011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100101010111110110100000001100011101011111011010000000110001110101111101101000000011000111010111110110100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 55600
ALLPIS = 62'b01110101011100010011101010000011111110001001001011000000101100;
XPCT = 39'b100000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 55900

pattern = 93; // 55900
LOAD0 = 112'b1010011011111011110111111111111101101110101011111011111100010010100000110000000000011111010000100000001110010101;
LOAD1 = 112'b0001001111110001100011000001110001010011101000010111100010001101000000111110010100101110011101110000110101011000;
LOAD2 = 112'b0101000111110000110111111110110101111111101100101011110000010100000001001110101100111110100011111111101010000011;
LOAD3 = 112'b0111100000010010101011001000011100010010011001010011101101000000000100101011001011110100111101001010111111010001;
UNLOAD[0] = 112'b1011011110110010110010010011100110100010101001100000110010000111010110100000001010101110001001110101000001111110;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100010111000111110100000100000010100101100001111101000001000000101001011011010100x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000110010110001111010000000000011001011000111101000000000001100101100001100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000010100011110100000000000110010110001111010000000000011001011000111101000000000001100101100011110100000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 56200
ALLPIS = 62'b01111010101110001001110101000001111111000100100101100000100110;
XPCT = 39'b000000000000000000000000000000101001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 56500

pattern = 94; // 56500
LOAD0 = 112'b0000010010111101111101111111111111101110111111011100010100111110001011111100000000001111101000100000001011001011;
LOAD1 = 112'b0110010011111100011000110000010011110100000101011110110000010010110100001111011010010110011011111001011011100001;
LOAD2 = 112'b0110000101010100001111110111010101100101010111001011111000111011010100101000001111001011101000111111111010100110;
LOAD3 = 112'b0110111100000010010101110100001010001101001001101000110110101000000010010001000111111110011110111001100101100001;
UNLOAD[0] = 112'b0000000000010101011100111010011001101000110010101011011011011111100000101000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000011001010000111101000000000001100101000011110100000000000110010100010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100010000001111010000000000011001010000111101000000000001100101000011110100000000000110010100001111010000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 56800
ALLPIS = 62'b01101101010111000100111010100000111111100010010010110000100011;
XPCT = 39'b100000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 57100

pattern = 95; // 57100
LOAD0 = 112'b1011011111011111110110111111111111111110110111110011010011001010011111000110101100000101110100100000001001100110;
LOAD1 = 112'b0101100100111101100110001100000101101011000010101111011000001001011010000111101101001011001101111100101100101011;
LOAD2 = 112'b0011010001111100000111111011100110110010101001100101111100011101101110011100001011110010111010001111101110101101;
LOAD3 = 112'b0111010000000001110110110010011000000110110011110100111110010011111001011010110010111101001111010010101111110100;
UNLOAD[0] = 112'b0000010011111101110001010011111000101111011010000101111101101111000011110100010110101011100010011101010000011111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101110111000001111101000100000001011001010000011111010001000000010110010111000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000001100100000011110100000000000110010000001111010000000000011001010000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100100100000111101000000000001100100000011110100000000000110010000001111010000000000011001000000111101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 57400
ALLPIS = 62'b01100110101011100010011101010000011111110001001001011000100001;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 57700

pattern = 96; // 57700
LOAD0 = 112'b0011111100111011100101110000000010110110100011001001100001011011101000011010010101101000001011111110001100011110;
LOAD1 = 112'b0010010010110001000000111010111110011101011110000110101111101000100111111100110000111110001011111111101110110100;
LOAD2 = 112'b0010110101011100001101110010001100011001101111010111000111100100000000001101110110111000001101000101000100000011;
LOAD3 = 112'b0110110000110001100100010110000000000011000101000101001101011010100100011011011111000111000010010011110111001010;
UNLOAD[0] = 112'b0000011011011111001101001100101001111100100001101101000110001110000100010110111000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001101000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000000000110011000001111010000000000011001100000111101000000000001100100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000100000010000011110100000000000110011000001111010000000000011001100000111101000000000001100110000011110100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 58000
ALLPIS = 62'b01101010011101110111110000111010101000110100010111010100101000;
XPCT = 39'b000000000000000000000000000000000000001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 58300

pattern = 97; // 58300
LOAD0 = 112'b1000010011001101111000111010000000011011000001100011001110111000011100001101000110110100000101011111001010001110;
LOAD1 = 112'b0110101110000100011000100110000111000111111111010111010011100101000110101111011100011110010000111010100101111111;
LOAD2 = 112'b0000010110100100001111010100000011110001111010010010110010111010010101101111111101101111000111010001010100000011;
LOAD3 = 112'b0100110010000001100010101011000000000001100010100010100110001101010110010111000001100000100000011001110011101111;
UNLOAD[0] = 112'b0111111000011001010111100100101101101101111110001111000011100111101001110000001000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b101000001011111110001100011111000011001000000000000000000000000000000000000000000000000000000000000000000000100x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111100010001111011010000101111110001000111101101000010111111000100011110001110110100000101111111000110001111101x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100101010110110100001011111100010001111011010000101111110001000111101101000010111111000100011110110100001011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 58600
ALLPIS = 62'b01110101001110111011111000011101010100011010001011101010101100;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 58900

pattern = 98; // 58900
LOAD0 = 112'b0010000000011110000010010100011110101110011011110000111001001110110010010000000010110011001001100001101101011001;
LOAD1 = 112'b0101010011110010100100010001010000101011100001000101001110111000101110001001010110110011101001101000011101001000;
LOAD2 = 112'b0110011000001010101101110001000101110100001001101110011101001100100010000011010101100110101100110000000101010001;
LOAD3 = 112'b0110000000110011000101110011110000000011110101010100011110111100001111001101101000110110110010110111001010111000;
UNLOAD[0] = 112'b0011111100000110001100111011100001110000011000110011001001110010010110100101010000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110100000101011111001010001111000001001110110100000101011111001010001111101101000001010111110010100011110000010x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111110001000111101101000010111111000100011110110100001011111100010001110011111011010000010101111100101000111110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110100111011010000101111110001000111101101000010111111000100011110110100001011111100010001111011010000101x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 59200
ALLPIS = 62'b01110000111010101010001100110100000010111001010010100001101110;
XPCT = 39'b000000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 59500

pattern = 99; // 59500
LOAD0 = 112'b0010001010001010100000011111110010101111100001100000010010011010100110110111000100110010101111001110110110110001;
LOAD1 = 112'b0001101100101111101011011100101110000001001110001100000000010110011010011010010011100101010101000001000000010111;
LOAD2 = 112'b0001111001011000100110101001111111010101011110111011111011000101000011101111001111100000110110011000010001000111;
LOAD3 = 112'b0000110011110011010110001111111100000010111111101111000010001100110111111101101011011100011011001000010010010110;
UNLOAD[0] = 112'b0000000000011110000010010100011110101110001100001110001011001101000111111000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001110000010110011001001100001101101011000101100110010011000011011010110010000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000011010101100101100100100100001101010110010110010010010000110101011000011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100110001011001001001000011010101100101100100100100001101010110010110010010010000110101011001011001001001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 59800
ALLPIS = 62'b01100010000000100010110110100000101001101000111110000100100111;
XPCT = 39'b000000000000000000000000000000000000000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 60100

pattern = 100; // 60100
LOAD0 = 112'b1100011000101010111101110111111110101000010111101110010111010111001100111110011111110000011100001001011011000111;
LOAD1 = 112'b0100100011011010011000101111110000011001111001101000100111000001000000010011110001001110001011010101101101101011;
LOAD2 = 112'b0010001001110001111011101100101101110100111001011100110100111110111001110100010001000000010000100010010100000110;
LOAD3 = 112'b0100100010111011101110010100100011111010110101000111110100110101101010100101101010101001001111110111111110000001;
UNLOAD[0] = 112'b1100001010000110000001001001101010011011001101001100110010100110000000100111010000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110010101111001110110110110001000000000000000000000000000000000000000000000000000000000000000000000000000000110x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011101111011001001100010111101110111101100100110001011110111011110110000011010011001010111100111011011011000100x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100111110110011000101111011101111011001001100010111101110111101100100110001011110111011110110010011000101111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 60400
ALLPIS = 62'b01101011011101100110101011101010111100000000001000010110101011;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 60700

pattern = 101; // 60700
LOAD0 = 112'b1100001001000101011110111011111111011100101011100110100010001111110110011110011111111010001110000100100101100011;
LOAD1 = 112'b0101001000110100100110001011111011000100111100110100010011100000100000001001111000100111000101101010110100100000;
LOAD2 = 112'b0101000100111000111101110110011010111010011110101110001010011111011100111110001100010100000100001000100101000001;
LOAD3 = 112'b0010100011100100011111001101001111000100101011001101000111101110111100110010110101010100100111111011111111000000;
UNLOAD[0] = 112'b0000011001011110111001011101011100110011100100100100101111011110011011010110100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000011000111110000011100001001011011000111111100000111000010010110110001110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010010101100011111100001110001001010110001111110000111000100101011000100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000110111011111000011100010010101100011111100001110001001010110001111110000111000100101011000111111000011100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 61000
ALLPIS = 62'b01100101101110110011010101110101011110000000000100001011101101;
XPCT = 39'b000000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 61300

pattern = 102; // 61300
LOAD0 = 112'b1111011111011001000010101111101101000001100010001001110110100001000100010010001010010100001100011100011110101111;
LOAD1 = 112'b0001101010011110101011111010000100111111000000010110000100110000110101011000000100001101001011000000010100111111;
LOAD2 = 112'b0000010111000001111000010011000010111110111101110010000000011111010101010000111001111101011100010110011001000111;
LOAD3 = 112'b0000100010101110011111001100111001110111100101001100010010101101000000000010000101101101010001101110001000101010;
UNLOAD[0] = 112'b0000001010101110011010001000111111011001101001100101001001000001010110110110100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001000011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001001010110001111110000111000100101011000111111000011100010010101100000010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111101011111100001110001001010110001111110000111000100101011000111111000011100010010101100011111100001110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 61600
ALLPIS = 62'b01111000101010101110011010000000000111110100010101010001101110;
XPCT = 39'b000000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 61900

pattern = 103; // 61900
LOAD0 = 112'b1111110110010100010000010011111100001100010001010010111011010010100010001000100101001011000110001110000111010110;
LOAD1 = 112'b0110011010100101101010111110101001011110110000011010010111011101001110101101000010010111100001100000001001010010;
LOAD2 = 112'b0100001011000110011100001001101001011111011101111001000000001011101110101110000010011111010111010101100110010011;
LOAD3 = 112'b0010100011110100011101010101010011110001110000010101000001100100100111011110001111101111101101101000101110001101;
UNLOAD[0] = 112'b1011111100011000010001100110000000000000100011111010111011010010001010000110010000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010100001100011100011110101111000111001000000000000000000000000000000000000000000000000000000000000000000000110x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111000111010110100101000110011100011101011010010100011001110001110101100011001001010000110001110001111010111010x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110101101001010001100111000111010110100101000110011100011101011010010100011001110001110101101001010001100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 62200
ALLPIS = 62'b01111100010101010111001101000000000011111010001010101000100111;
XPCT = 39'b000000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 62500

pattern = 104; // 62500
LOAD0 = 112'b0111111011110110010101010100111100001110101011101100111100110011111001011010010011001100101000011001001111110111;
LOAD1 = 112'b0111110110111010010010110111010101101111000110000011100110000110101010000000111011011111110011100111101001100100;
LOAD2 = 112'b0110110000101100010000100100000000100100111100100001010111010011010000010100110010011011111001110001001100100111;
LOAD3 = 112'b0010001010101010101010001100101001110111111101001111101101000000100011111011111110011100010110001000010101000000;
UNLOAD[0] = 112'b0101100010010100010000010011111100001100001110101110101000101000000000000100111000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001011011101001011000110001110000111010111010010110001100011100001110101110000111x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011100011101011010010100011001110001110101101001010001100111000111010100010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111111010100101000110011100011101011010010100011001110001110101101001010001100111000111010110100101000110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 62800
ALLPIS = 62'b01100100010111011100010110011010101001001001010010000000100011;
XPCT = 39'b000000000000000000000000000000000000110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 63100

pattern = 105; // 63100
LOAD0 = 112'b1001001111011111101110000011011000001100110101101010011110011010111100100000011101100101010100001100100011111011;
LOAD1 = 112'b0111010111101100101110001101111010111110100011010001110110010010010101000100001100111011101000100010100100010101;
LOAD2 = 112'b0011011000010110111100010110010111100110001101101100011010111010100000010100011000100111111010011100000010011110;
LOAD3 = 112'b0111101010100100010111101000100000011111111010000010111110001111000101011101111111001110001011000100001010100000;
UNLOAD[0] = 112'b0000011110111001101101000100100110000001000111011110000110111101001100101000000010001011101110001011001101010101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b001100101000011001001111110111000000001011001100101000011001001111110110110011001010000110010011111101111000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110010011111010110011010100011001001111101011001101010001100100111110101000001100110010100001100100111111011011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000001100110101000110010011111010110011010100011001001111101011001101010001100100111110101100110101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 63400
ALLPIS = 62'b01110010001011101110001011001101010100100100101001000000101001;
XPCT = 39'b000000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 63700

pattern = 106; // 63700
LOAD0 = 112'b1000101000111101011010011101101001000110111010101011001111001100011110011010010110110001101010000110010001111100;
LOAD1 = 112'b0101110101111011101011100011011011011010110001101000111011001001001010100010000110011101110100010001010001111001;
LOAD2 = 112'b0001101100001011110110001011001111110011000101110110001101001101011000011011011110001000111110110111000000100001;
LOAD3 = 112'b0111000110010110101010110010110010011100000100110111111100110001011010001110111111100111000101100010000101010000;
UNLOAD[0] = 112'b0000011111011111101110000011011000001100000001100111101110101101110001110100100001000101110111000101100110101011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000100111011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011001001111101011001101010001100100111110101100110101000110010011111001000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110100110110011010100011001001111101011001101010001100100111110101100110101000110010011111010110011010100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 64000
ALLPIS = 62'b01111001000101110111000101100110101010010010010100100000100100;
XPCT = 39'b100000000000000000000000000001100011101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 64300

pattern = 107; // 64300
LOAD0 = 112'b1100001110110100100001101110100101000000011110000010000110111100100111011011100110110010111110111101001000100010;
LOAD1 = 112'b0001100101001111011000100000000111101101000110011010111010101110101000001111111011110010011011111101100101011100;
LOAD2 = 112'b0010000011011000010101101101100100011010010001011110100011110110010111001010011101011010010010101001110000001011;
LOAD3 = 112'b0010001100100100101011010011000001001100110011101100110100011110110101111100000000110100100000100010110101100010;
UNLOAD[0] = 112'b0000001000111101011010011101101001000110101111001110010001010001111110101000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001100100111111101100110101000110010011111110110011010100011001001111100011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000110010111011001101010001100100111111101100110101000110010011111110110011010100011001001111111011001101010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 64600
ALLPIS = 62'b01110110111111001100010010001001111101111101011101000100101010;
XPCT = 39'b100000000000000000000000000000000001000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 64900

pattern = 108; // 64900
LOAD0 = 112'b0101011001011101100110101011110110000000001100011000100010000100111011110001110010110010010100010000100100001101;
LOAD1 = 112'b0100100001000000010100010000111110110011111111100001011000010111010001111001000111100101100100001011011101101010;
LOAD2 = 112'b0011110100110001100010111000111111111100011110010101101101011101110111001111100101101011111001101110011100010011;
LOAD3 = 112'b0011100010100001100100101001100100101001011110011010100101111010101010000101011111011101010010000010101101111011;
UNLOAD[0] = 112'b1000101010110100100001101110100101000000101001101100001001011010110111110111110011011111100110001001000100111110;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110010111110111101001000100011100000001110110010111110111101001000100011101100101111101111010010001000110010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111010000010001101100011111011101000001000110110001111101110100000100010000011011001011111011110100100010001110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000000011011000111110111010000010001101100011111011101000001000110110001111101110100000100011011000111110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 65200
ALLPIS = 62'b01110001000010010001111001111110010110001010111001110110100101;
XPCT = 39'b000111111100001011000010111010001110100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 65500

pattern = 109; // 65500
LOAD0 = 112'b1001011100101011110001011101101110010000000110000110010001000011011101111000010001011010001010101000010010000101;
LOAD1 = 112'b0111001000010000000101000100001011011100000100010001110101101100001100001100101000000000011110001101111110001101;
LOAD2 = 112'b0101111010011000111011101001010010110111100000010111100110110100101010111101111101011010111110001011110111000010;
LOAD3 = 112'b0110110111000011100010100100110110010000101111001101010010111101010101000010101111101110101001000001010110111101;
UNLOAD[0] = 112'b0000011011110001101000010000000110001111101100010010100100011000111000011000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100001010000110101100001010010000101000011010110000101001000010100001100011100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000110100001011000010100100001010000110101100001010010000101000011010110000101001000010100001101011000010100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 65800
ALLPIS = 62'b01111000100001001000111100111111001011000101011100111011101010;
XPCT = 39'b100000000000000000000000000000000001111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 66100

pattern = 110; // 66100
LOAD0 = 112'b1110111111111110011001010110110101100111100000001000101001111001000110100001001101000110001110011010000001011110;
LOAD1 = 112'b0111001010010111100011001001110001111110010001110100010011000101110011000010001011101101011000011101010010001111;
LOAD2 = 112'b0100001000010001101001101111100000111000011111100111110100001110001100000110010101101111110010100110111101100001;
LOAD3 = 112'b0000001000111101011000111001010110111100000011010011100101001001000000011010001000110000010110110011011100010100;
UNLOAD[0] = 112'b0000011010010000010011001101011010010000010011001100101100101010010111100100100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010100000000001111000110111110001011011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010000101000010010110000101001000010100001001011000010100100001010000100001100010001000111010110110000110000110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100111000100101100001010010000101000010010110000101001000010100001001011000010100100001010000100101100001010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 66400
ALLPIS = 62'b01100110001101010011101110100101001101010110111001001001101101;
XPCT = 39'b000000000000000000000000000000000001110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 66700

pattern = 111; // 66700
LOAD0 = 112'b0101001010010111000011100000011111000111110000010010010100111100100011010011000110100011000111101101000000101100;
LOAD1 = 112'b0011110010100101011000110010010011111011101100111011001100110110101101100100010100110110111101011011111010010010;
LOAD2 = 112'b0010000100001001110100110001001011110001000101100010001011110000000010110010001101011110111100111001101111011000;
LOAD3 = 112'b0001101011110001001010011010011011101011101010010001010010100110001011101101000100011000001011011001101110001010;
UNLOAD[0] = 112'b0000011110101100011100000010100000010001110100000101011110000110010111000101010011000110101001110111010010100111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110100000101111010001000111011010000010111101000100011101101000001011101000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100000000010100010001110110100000101111010001000111011010000010111101000100011101101000001011110100010001110x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 67000
ALLPIS = 62'b01110011000110101001110111010010100110101011011100100100100110;
XPCT = 39'b000000000000000000000000000000000000000;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 67300

pattern = 112; // 67300
LOAD0 = 112'b0111110000110100001110101001101001101010000001000000101000011011100001011111110110111000101000001000100100001010;
LOAD1 = 112'b0010000100111000110100010100010111100000001000110011000001010001011011101100110010100111111111011000110001111100;
LOAD2 = 112'b0111101011100111101000110011110011101101110111011100111000001101011010000101101101101111110010011010011011100011;
LOAD3 = 112'b0111010111111100000001011011001001111010110000001100100100001001100101000001111100110111010000100111110011001010;
UNLOAD[0] = 112'b0000001010010111000011100000011111000111101110100101011110001110010001011000000001100011010100111011101001010011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011010000010111101000100011101101000001011110100010001110110100000101100010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000111110011010001000111011010000010111101000100011101101000001011110100010001110110100000101111010001000111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 67600
ALLPIS = 62'b01110011111110100011001011010011111011100001111001000110100011;
XPCT = 39'b100000000000000000000000000100011110011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 67900

pattern = 113; // 67900
LOAD0 = 112'b0001100000000100000010101001010101111000001110101011110100111000110100101000011010110110011111111010011110011011;
LOAD1 = 112'b0100011001011111001111011101110000110101111010110111000111100010100000101000100001101111011110011001010111001010;
LOAD2 = 112'b0111001110110001010000111100011010010001001011011101000111010010010010111001011101100110100001110010110110101101;
LOAD3 = 112'b0010111110001000100100001011100000111110011001000011001111111110000010101101100001100010100001101100010111001101;
UNLOAD[0] = 112'b0000010000000100000010100001101110000101010100101100000111101111101100010100000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b011001010011111111101100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b010001010000101101110010100001000101000010110111001010000100010100001000000000100011001100000101000101101110110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000011011100101000010001010000101101110010100001000101000010110111001010000100010100001011011100101000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 68200
ALLPIS = 62'b01100011100010100110010101010011010101000100101011110111100001;
XPCT = 39'b100000000000000000000000000000000000110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 68500

pattern = 114; // 68500
LOAD0 = 112'b0010110101101110110001011100010110110101100111001011111011001101101100001110000101011011001111111101001111001111;
LOAD1 = 112'b0011000110010111110011110111011101001111011101011011100011110001010000010100010000110111101111001100101000000011;
LOAD2 = 112'b0111100111011110011001011000111101001010100110100101110100100011000111011010101111011100101000011100111101101001;
LOAD3 = 112'b0111011000100100000010100101100100010111001101100000110111011111010001010111110000110101010000100110001011100000;
UNLOAD[0] = 112'b0001100000000100000010101001010101111000000001010101000110101001011111011000000001110001010011001010101001101010;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010000110111101111001100101010000110101010110110011111111010011110011010101101100111111110100111100110110010010x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110100111001100101101001111111010011100110010110100111111101001110011010001011101011011100011110001010000010100x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010010101101011010011111110100111001100101101001111111010011100110010110100111111101001110011001011010011111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 68800
ALLPIS = 62'b01100001110001010011001010101001101010100010010101111011101000;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 69100

pattern = 115; // 69100
LOAD0 = 112'b1110011001100111011100100110011010011011010011110011111101001111001101000000110110101100100111111110101011100111;
LOAD1 = 112'b0010110001100101011100111101110100110110001100000101110001111000100000000010000000110011111101001110011110100111;
LOAD2 = 112'b0011110011101100100100101100001110100101010011010010111010010101100011100001001011110111001010010111001111011010;
LOAD3 = 112'b0111111110010100000100011110000110110011000110111100100110001110011010001011011000011000101000011011000101110011;
UNLOAD[0] = 112'b0000010010011100101111101100110110110000011100001110111110110001100100110110011000111000101001100101010100110101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001001001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111010011100111010110100111111101001110011101011010011111110100111001100010100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100100110101101001111111010011100111010110100111111101001110011101011010011111110100111001110101101001111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 69400
ALLPIS = 62'b01100000111000101001100101010100110101010001001010111101101100;
XPCT = 39'b100000000000000000000000000000000001001;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 69700

pattern = 116; // 69700
LOAD0 = 112'b1110001010100110101110010000011001000000101001111101111110100101100110101000000111010101010011011111011001110010;
LOAD1 = 112'b0100101100011011010111001111011101011011010111010110111000111100010100000101000100001101111011110011001000110100;
LOAD2 = 112'b0101111001110110010010010110000111010010101010101001101101011010110001101100111110111101110010110101100011110100;
LOAD3 = 112'b0111100101010010010000010101001110000011110000011001000101011111101110100101101100001100010100001101100010111001;
UNLOAD[0] = 112'b0000011111001000111101010000011010100000000100101011110100111001001101001000000000011100010100110010101010011011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000110111000000000000000000000000000000000000000000000000000000000000000001000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111101001110011101011010011111110100111001110101101001111111010011100100001000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110010111010110100111111101001110011101011010011111110100111001110101101001111111010011100111010110100111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 70000
ALLPIS = 62'b01100000011100010100110010101010011010101000100101011110101110;
XPCT = 39'b100000000000000000000000000100111001111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 70300

pattern = 117; // 70300
LOAD0 = 112'b0111010010000110011011001111101001101110010100111110111111010001110011010001101111101001101001011111100100111011;
LOAD1 = 112'b0001001011000100110101110011110011110100101011101011011100011110001010000010100010000110111101111001100101110100;
LOAD2 = 112'b0111110100110011000001001011001011101001010100010100110110111001011100101111011011101111011100111101001000111111;
LOAD3 = 112'b0100010101001010010000001000100011101001111000011100100010001111110110110111110111000101011000100010111001011111;
UNLOAD[0] = 112'b0000011110100110101110010000011001000000100000011010101011111111100001001000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001011000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111110100111001110101101001111111010011100111010110100111111101001110000000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100101010011101011010011111110100111001110101101001111111010011100111010110100111111101001110011101011010011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 70600
ALLPIS = 62'b01100000001110001010011001010101001101010100010010101111101111;
XPCT = 39'b100000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 70900

pattern = 118; // 70900
LOAD0 = 112'b0001111100010001101010010011010111011110001001010110111110110001010001110011011010011100111111100001111110000010;
LOAD1 = 112'b0110001000100000101111000110001001110111000011110011001001000111000000011101100001111111110101001011111101001100;
LOAD2 = 112'b0001101011000000100110001101101110000111011001101111100010001010010101111011001101000110101110011010010010011011;
LOAD3 = 112'b0100100000011010111100010010000101110011111000001011001100111101001011000010000100000100000111010000101111100100;
UNLOAD[0] = 112'b1110110010000110011011001111101001101110001010100011100111011111011100001000000000000000000000000000000000000000;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010001000011011110111100110010000000011111101001101001011111100100111011111010011010010111111001001110110000100x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111111010011101111010110100111111101001110111101011010011111110100111010000010101110101101110001111000101000001x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011110101101001111111010011101111010110100111111101001110111101011010011111110100111011110101101001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 71200
ALLPIS = 62'b01111010011010110010111100010000001110011110011110000011101111;
XPCT = 39'b000000000000000000000000000000000000101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 71500

pattern = 119; // 71500
LOAD0 = 112'b0001111000110011010110110011101000000001000111101100111110000001000000100010111000100111010100101110110011011100;
LOAD1 = 112'b0111010010111001101001101001111111100011101011100011000011101000101001010001001100000011011110011001110000000101;
LOAD2 = 112'b0010000000111101101101101110011101101000011100010010110010000100110101010100000100101100110011110010110100100011;
LOAD3 = 112'b0110101001010101111010111111000010110110111100000001111011001100010101111010011101000101000001111011100000111000;
UNLOAD[0] = 112'b0000011111111010111101110100000011101101000101111000100101001101000001110111100000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001110101010011100111111100001111110000010100111001111111000011111100000110000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000011111000000100111011111100001111100000010011101111110000111110000010011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100011001001110111111000011111000000100111011111100001111100000010011101111110000111110000001001110111111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 71800
ALLPIS = 62'b01100111010000101110101110110010101111111011011000010101101111;
XPCT = 39'b000000000000000000000000000000000000101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 72100

pattern = 120; // 72100
LOAD0 = 112'b1010010000110111001000101011100111110110101110110011111110111010000100011100011101111001100001011001010001110011;
LOAD1 = 112'b0101000100111111011000000010101100100001101011001111000110111110011001110110011110111101001110111101110110001001;
LOAD2 = 112'b0001101101001011110000011111011001110111111101101100101100000110101101110100101011110111010000111000101101011111;
LOAD3 = 112'b0011011000101111001001111001110001010100011110000101100000110100101110100000110001000100100000110110010111010111;
UNLOAD[0] = 112'b0000011100000011101100101011011110010001110000100011011110011111000111001000000011101000010111010111011001010111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b100111010100101110110011011101101100000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011101101101110001001101010001110110110111000100110101000111011011011101010100010011101010010111011001101110000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100101010100010011010100011101101101110001001101010001110110110111000100110101000111011011011100010011010100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 72400
ALLPIS = 62'b01111001110101100000100111100011111111001001111011011110101111;
XPCT = 39'b000000000000000000000000000000000001100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 72700

pattern = 121; // 72700
LOAD0 = 112'b1110011011001110101010001101100110111011110000001101111111001100100100001000010110111110110000011100100100111000;
LOAD1 = 112'b0111010001001111110110000000100110001101010101100111101011011101101100011011001111011110000111011110111000000111;
LOAD2 = 112'b0001111010100001011000001111101100111011111111110110000110010011010010110001010110111101110100011110001011010011;
LOAD3 = 112'b0111000111110110111100011100111100100110001001000110100100110010010111010011001000110010110001010111000011101011;
UNLOAD[0] = 112'b0000010010111011001111111011101000010001000110011011110011000101010111010100100100111010110000010011110001111111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110010100111001011110110000111001010011100101111011000011100101001110001000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000000101110111101100001110010100111001011110110000111001010011100101111011000011100101001110010111101100001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 73000
ALLPIS = 62'b01111100111010110000010011110001111111100100111101101111100111;
XPCT = 39'b100000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 73300

pattern = 122; // 73300
LOAD0 = 112'b0101011101001000111110110100110100101011101010011011011110111100011010001110111110110101010011010000011110000011;
LOAD1 = 112'b0101001100000010011111111000110110011011010100011101010110100101101011000011011111010011110010011010010010001010;
LOAD2 = 112'b0110001000001100101010101111111101111111001101011110000100001101101010011111000011010011000000010011110010100111;
LOAD3 = 112'b0010110110101111011110111000001110011000000100100100111101101011111111110010111011011110011010111000010110111111;
UNLOAD[0] = 112'b0000011010111100100110101110011010110011000001100111001001101101011000101000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111001010011101101111011000011100101001110110111101100001110010100111000000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100100000011011110110000111001010011101101111011000011100101001110110111101100001110010100111011011110110000x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 73600
ALLPIS = 62'b01110100000000101111111001000010010111000110001001100011101011;
XPCT = 39'b100000000000000000000000000000000000110;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 73900

pattern = 123; // 73900
LOAD0 = 112'b0011100010001001010111011010011110001101101101110111101111011111011101000010100111011011101001011000000111000010;
LOAD1 = 112'b0111010011000000000111111110001111010101101010001110101011010010110101100001101111101001111001001101001010001110;
LOAD2 = 112'b0111000100000110101001000111110110111111000101101111010011001010101111011000101100110101110000000100101100101101;
LOAD3 = 112'b0110010011110101111111001100010011001100000110010010001110111101101111011001011101101111001101011100001011011111;
UNLOAD[0] = 112'b0000011010101001101101111011110001101000000101110100000010100110101001000111000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b110101010011010000011110000011000011000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100000111000001101101101001110000011100000110110110100111000001110000010011011011010101001101000001111000001110x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000100010011011011010011100000111000001101101101001110000011100000110110110100111000001110000011011011010011x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 74200
ALLPIS = 62'b01111010000000010111111100100001001011100011000100110001100101;
XPCT = 39'b000000000000000000000000000000000000111;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 74500

pattern = 124; // 74500
LOAD0 = 112'b0010101110001111000000000111001001100000110101100100010010110110000110111110111010000110111111000010001111111111;
LOAD1 = 112'b0001001100100001100011100111010011111010101011101001110010100011010111101110001111001000011101010011101010001010;
LOAD2 = 112'b0101010111011111001010000011110100111100010011110011110100110101000100111100110101110101000001010101011011011100;
LOAD3 = 112'b0010101011101100001011100000001001100001000011001100011010001100010011110111110001110000100100111101110010100101;
UNLOAD[0] = 112'b0000000010001001010111011010011110001101011001110011000101111000110001101000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b011011101001011000000111000011000000001000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110000011100001110110110100111000001110000111011011010011100000111000000000011101101110100101100000011100001111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100100000011101101101001110000011100001110110110100111000001110000111011011010011100000111000011101101101001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 74800
ALLPIS = 62'b01100111011101111100001110101010001101000101110101001100100010;
XPCT = 39'b000000000000000000000000000000000000010;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 75100

pattern = 125; // 75100
LOAD0 = 112'b0000011011010011101000000001110001101000011010101000001011011011000011010111011101000011011111110001000011111111;
LOAD1 = 112'b0000010011001010011000111001111011111001110101110100111001010001101011110111000111100100001110101001110100001000;
LOAD2 = 112'b0110101011101111110101000001111100011110001000101001101010011110110000001010011001011001010000010101010110110111;
LOAD3 = 112'b0111111010111110000101010000010000111000100000100111001101000110001001011011111000111000010010011110111001010010;
UNLOAD[0] = 112'b0000001011010110010001001011011000011011010111111001110110011101100010110111001011101110111110000111010101000111;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b000100011111110100001011111100010001111111010000101111110001000111111101000100000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000011110001000010111111000100011111110100001011111100010001111111010000101111110001000111111101000010111111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 75400
ALLPIS = 62'b01110011101110111110000111010101000110100010111010100110100001;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 75700

pattern = 126; // 75700
LOAD0 = 112'b1100011010111000111010000000101100101100001101001010000101101110100001101000000110100010101111111000101001111101;
LOAD1 = 112'b0110000100110000100110001110011101101100111010011010011100101000110101110011100011110010100111010100111010101011;
LOAD2 = 112'b0011010101110111111010100000111110001111000110010100010101011011011100011011011110010111010100000101000101101101;
LOAD3 = 112'b0111110111110001010011011000011000000100010100010110110110011011000000101101111100011100001001001111011100101001;
UNLOAD[0] = 112'b0000011001101010100000101101101100001101010010101000110110000010100111000111100001110111011111000011101010100011;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101111000000000000000000000000000000000000000000000000000000000000000000000010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b100010001111111010000101111110001000111111101000010111111000100011111100010000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000010111110100001011111100010001111111010000101111110001000111111101000010111111000100011111110100001011111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 76000
ALLPIS = 62'b01101001110111011111000011101010100011010001011101010011100000;
XPCT = 39'b100000000000000000000000000000000001101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 76300

pattern = 127; // 76300
LOAD0 = 112'b1110011111011101010111000000000111001110000110100011000010110101010000110000100011010010010111111100011000111111;
LOAD1 = 112'b0011100001001110001001100011101100101011111101011101001110010100111010110101110001111001000011101010011110100111;
LOAD2 = 112'b0101101010111011011101010000011111000111100011001010101010101001101110001111101011100001110101010001000001011101;
LOAD3 = 112'b0110110110001101001001001100000000001110001010001010011001000101100000110110111110001110000100100111101110010100;
UNLOAD[0] = 112'b0000011001101011001101111101010110101010000101000000101101011000001111101000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000001101011000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b110001000111111101000010111111000100011111110100001011111100010001111100011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001000111110011010000101111110001000111111101000010111111000100011111110100001011111100010001111111010000101111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 76600
ALLPIS = 62'b01110100111011101111100001110101010001101000101110101001100000;
XPCT = 39'b100000000000000000000000000000000001011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 76900

pattern = 128; // 76900
LOAD0 = 112'b0011100110111010100111111111011100100011101000101001110100010101111110110100101001001111110100001110010010011001;
LOAD1 = 112'b0010100101010000100101000001101011011010101011011010000011010101001010001111111110111010001011000110001100101000;
LOAD2 = 112'b0111111100000001101101100100100101110100100100010011011101001110011010010100110001000001110000001011110001101110;
LOAD3 = 112'b0110011001011000011010001011011111011011000010111011111100001010101010100000110101111011011001001110110101111010;
UNLOAD[0] = 112'b0000011110001111101010010111100011001010110111101001100111000011000101110100111000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b010010010111111100011000111111000101000000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b111000100011110110100001011111100010001111011010000101111110001000111110011101101001001011111110001100011111011x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000100110110001101000010111111000100011110110100001011111100010001111011010000101111110001000111101101000010111x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 77200
ALLPIS = 62'b01110000011100101000011011001010110101101010110010100011100010;
XPCT = 39'b000000000000000000000000000000000000011;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 77500

pattern = 129; // 77500
LOAD0 = 112'b0000111000011101011001111111111011001000110100011010111010001011111111011011100000100111111010100111000101001100;
LOAD1 = 112'b0100101001010110001001010000010111110000110101101101000001101010100101000111111111011101000101100011000100101000;
LOAD2 = 112'b0011111110000000011110110010010010111010010001001001011110100011101101000111000100010000011100000010101100011111;
LOAD3 = 112'b0111001001101101001101000101101011101101100100011101111110100101000101110000011010111101101100100111011010111101;
UNLOAD[0] = 112'b0011100010100010100111010001010111111011111010101111111110010101010111000100111000001110010100001101100101011010;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b111111011101000101100011000110101011000001111111110101100111100101100011011110111001011000010011111100101010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011100101001100010011111010001110010100110001001111101000111001010011001000110101101101000001101010100101000111x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000010001011000100111110100011100101001100010011111010001110010100110001001111101000111001010011000100111110100x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 77800
ALLPIS = 62'b01111000001110010100001101100101011010110101011001010001101001;
XPCT = 39'b000000000000000000000000000000000000101;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 78100

pattern = 130; // 78100
LOAD0 = 112'b0111011001110001000001010000100001010111110010101110101001010011000001001000011001011100001001101101111000111101;
LOAD1 = 112'b0101101111000111100111010101101000110010110001001100100011100000111000101100000011010100101001110111101110000111;
LOAD2 = 112'b0010000011000001001010011101101000101001101100110101000010001011111000100000001000000100110111001011011010101111;
LOAD3 = 112'b0011110111100001111100011001111010101001110100110101010011101000001000111000111000100101101111011101011000100100;
UNLOAD[0] = 112'b0000011000101011100101000011010001010101110000111111100100110000001101101000000100000111001010000110110010101101;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000101110100000000000000000000000000000000000000000000000000000000000000000001010000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b001110010100110001001111101000111001010011000100111110100011100101001101011000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b000000001101100010011111010001110010100110001001111101000111001010011000100111110100011100101001100010011111010x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 78400
ALLPIS = 62'b01101100011011100010011101111000011000110000011110001011101110;
XPCT = 39'b100000000000000000000000000000000000100;
MASK = 39'b111111111111111111111111111111111111111;
#0 ->capture_hclk;
#300; // 78700

lastpattern = 1;
LOAD0 = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
LOAD1 = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
LOAD2 = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
LOAD3 = 112'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
UNLOAD[0] = 112'b0000011101111111110011001000001011001000001010111011110101011110100111001000000000000000000000000000000000000001;
UNLMSK[0] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
UNLOAD[1] = 112'b000000000000000000000000000000000110100000000000000000000000000000000000000000000000000000000000000000000000000x;
UNLMSK[1] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[2] = 112'b011011100011110010111000100101101110001111001011100010010110111000111100000000000000000000000000000000000000000x;
UNLMSK[2] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
UNLOAD[3] = 112'b001100111100000101110001001011011100011110010111000100101101110001111001011100010010110111000111100101110001001x;
UNLMSK[3] = 112'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110;
#0 ->load_unload;
#load_delay; // 79000
      $display("// %t : Simulation of %0d patterns completed with %0d errors\n", $time, pattern+1, nofails);
      if (verbose >=2) $finish(2);
      /* else */ $finish(0);
   end
endmodule
