module ctrl;

// 0in set_cdc_reconvergence_depth 10

// 0in set_cdc_clock hclk -period 50

endmodule

